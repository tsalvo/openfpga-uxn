-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 59
entity nip2_0CLK_15c648e1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_15c648e1;
architecture arch of nip2_0CLK_15c648e1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2307_c6_98c3]
signal BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2307_c1_a907]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2307_c2_96b3]
signal result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2307_c2_96b3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2307_c2_96b3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2307_c2_96b3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2307_c2_96b3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2307_c2_96b3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l2307_c2_96b3]
signal t16_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l2308_c3_8e53[uxn_opcodes_h_l2308_c3_8e53]
signal printf_uxn_opcodes_h_l2308_c3_8e53_uxn_opcodes_h_l2308_c3_8e53_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2312_c11_f7d9]
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2312_c7_d7c4]
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2312_c7_d7c4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2312_c7_d7c4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2312_c7_d7c4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2312_c7_d7c4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2312_c7_d7c4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l2312_c7_d7c4]
signal t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2315_c11_0d39]
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2315_c7_37fa]
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c7_37fa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c7_37fa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2315_c7_37fa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2315_c7_37fa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c7_37fa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l2315_c7_37fa]
signal t16_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2317_c3_994b]
signal CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2320_c11_0f80]
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2320_c7_ca68]
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2320_c7_ca68]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2320_c7_ca68]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2320_c7_ca68]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2320_c7_ca68]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2320_c7_ca68]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l2320_c7_ca68]
signal t16_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2323_c11_627e]
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2323_c7_4765]
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2323_c7_4765]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2323_c7_4765]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2323_c7_4765]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2323_c7_4765]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2323_c7_4765]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l2323_c7_4765]
signal t16_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2324_c3_c7d9]
signal BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2326_c30_4259]
signal sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2331_c11_89a6]
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2331_c7_e873]
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2331_c7_e873]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2331_c7_e873]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2331_c7_e873]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2331_c7_e873]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(3 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l2334_c31_09f7]
signal CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2336_c11_b0c5]
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2336_c7_77a2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2336_c7_77a2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_25e8( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3
BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_left,
BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_right,
BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3
result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3
result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3
result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3
result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output);

-- t16_MUX_uxn_opcodes_h_l2307_c2_96b3
t16_MUX_uxn_opcodes_h_l2307_c2_96b3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2307_c2_96b3_cond,
t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue,
t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse,
t16_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output);

-- printf_uxn_opcodes_h_l2308_c3_8e53_uxn_opcodes_h_l2308_c3_8e53
printf_uxn_opcodes_h_l2308_c3_8e53_uxn_opcodes_h_l2308_c3_8e53 : entity work.printf_uxn_opcodes_h_l2308_c3_8e53_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2308_c3_8e53_uxn_opcodes_h_l2308_c3_8e53_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_left,
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_right,
BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4
result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4
result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output);

-- t16_MUX_uxn_opcodes_h_l2312_c7_d7c4
t16_MUX_uxn_opcodes_h_l2312_c7_d7c4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond,
t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue,
t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse,
t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_left,
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_right,
BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_cond,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output);

-- t16_MUX_uxn_opcodes_h_l2315_c7_37fa
t16_MUX_uxn_opcodes_h_l2315_c7_37fa : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2315_c7_37fa_cond,
t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue,
t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse,
t16_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2317_c3_994b
CONST_SL_8_uxn_opcodes_h_l2317_c3_994b : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_x,
CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_left,
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_right,
BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_cond,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68
result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68
result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output);

-- t16_MUX_uxn_opcodes_h_l2320_c7_ca68
t16_MUX_uxn_opcodes_h_l2320_c7_ca68 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2320_c7_ca68_cond,
t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue,
t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse,
t16_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_left,
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_right,
BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_cond,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_return_output);

-- t16_MUX_uxn_opcodes_h_l2323_c7_4765
t16_MUX_uxn_opcodes_h_l2323_c7_4765 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2323_c7_4765_cond,
t16_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue,
t16_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse,
t16_MUX_uxn_opcodes_h_l2323_c7_4765_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9
BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_left,
BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_right,
BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2326_c30_4259
sp_relative_shift_uxn_opcodes_h_l2326_c30_4259 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_ins,
sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_x,
sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_y,
sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_left,
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_right,
BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_cond,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873
result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873
result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_return_output);

-- CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7
CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_x,
CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_left,
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_right,
BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
 t16_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output,
 t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output,
 t16_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output,
 CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output,
 t16_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_return_output,
 t16_MUX_uxn_opcodes_h_l2323_c7_4765_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_return_output,
 sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_return_output,
 CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iffalse : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_9c80 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2308_c3_8e53_uxn_opcodes_h_l2308_c3_8e53_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_6df0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_ee1a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2321_c3_d079 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2328_c3_d7c7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2329_c21_45c5_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2333_c3_0823 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_e873_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2334_c21_0949_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_f119_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2323_l2320_l2315_l2312_l2307_DUPLICATE_044d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_9c90_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2324_DUPLICATE_9d92_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2341_l2303_DUPLICATE_bafb_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2321_c3_d079 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2321_c3_d079;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2328_c3_d7c7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2328_c3_d7c7;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_9c80 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2309_c3_9c80;
     VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_6df0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2313_c3_6df0;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2333_c3_0823 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2333_c3_0823;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_ee1a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2318_c3_ee1a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_left := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_x := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea_return_output := result.is_opc_done;

     -- CONST_SR_8[uxn_opcodes_h_l2334_c31_09f7] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_x <= VAR_CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_return_output := CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2315_c11_0d39] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_left;
     BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output := BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2336_c11_b0c5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2320_c11_0f80] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_left;
     BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output := BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2307_c6_98c3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_9c90 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_9c90_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2312_c11_f7d9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_f119 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_f119_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2323_l2320_l2315_l2312_l2307_DUPLICATE_044d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2323_l2320_l2315_l2312_l2307_DUPLICATE_044d_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2331_c11_89a6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2324_DUPLICATE_9d92 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2324_DUPLICATE_9d92_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- sp_relative_shift[uxn_opcodes_h_l2326_c30_4259] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_ins;
     sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_x;
     sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_return_output := sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b_return_output := result.is_stack_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2331_c7_e873] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_e873_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2323_c11_627e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2307_c6_98c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2312_c11_f7d9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2315_c11_0d39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2320_c11_0f80_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2323_c11_627e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2331_c11_89a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2336_c11_b0c5_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2324_DUPLICATE_9d92_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2316_l2324_DUPLICATE_9d92_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2323_l2320_l2315_l2312_l2307_DUPLICATE_044d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2323_l2320_l2315_l2312_l2307_DUPLICATE_044d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2323_l2320_l2315_l2312_l2307_DUPLICATE_044d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2323_l2320_l2315_l2312_l2307_DUPLICATE_044d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2323_l2320_l2315_l2312_l2307_DUPLICATE_044d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2331_l2323_l2320_l2315_l2312_l2336_DUPLICATE_39ea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_9c90_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_9c90_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_9c90_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_9c90_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_9c90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_l2336_DUPLICATE_0c1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_f119_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_f119_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_f119_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_f119_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2331_l2320_l2315_l2312_l2307_DUPLICATE_f119_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2331_c7_e873_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2326_c30_4259_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2307_c1_a907] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2323_c7_4765] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2317_c3_994b] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_return_output := CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2334_c21_0949] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2334_c21_0949_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l2334_c31_09f7_return_output);

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2331_c7_e873] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2331_c7_e873] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2336_c7_77a2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2324_c3_c7d9] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_left;
     BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_return_output := BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2336_c7_77a2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2334_c21_0949_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2317_c3_994b_return_output;
     VAR_printf_uxn_opcodes_h_l2308_c3_8e53_uxn_opcodes_h_l2308_c3_8e53_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2307_c1_a907_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2336_c7_77a2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2320_c7_ca68] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2323_c7_4765] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2323_c7_4765] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2331_c7_e873] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2331_c7_e873] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;

     -- t16_MUX[uxn_opcodes_h_l2323_c7_4765] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2323_c7_4765_cond <= VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_cond;
     t16_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue;
     t16_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_return_output := t16_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2331_c7_e873] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_return_output := result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2329_c21_45c5] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2329_c21_45c5_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l2324_c3_c7d9_return_output);

     -- printf_uxn_opcodes_h_l2308_c3_8e53[uxn_opcodes_h_l2308_c3_8e53] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2308_c3_8e53_uxn_opcodes_h_l2308_c3_8e53_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2308_c3_8e53_uxn_opcodes_h_l2308_c3_8e53_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2329_c21_45c5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2331_c7_e873_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2320_c7_ca68] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2323_c7_4765] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_return_output := result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2315_c7_37fa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2320_c7_ca68] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2323_c7_4765] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2323_c7_4765] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;

     -- t16_MUX[uxn_opcodes_h_l2320_c7_ca68] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2320_c7_ca68_cond <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_cond;
     t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue;
     t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output := t16_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2323_c7_4765_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2320_c7_ca68] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2315_c7_37fa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2320_c7_ca68] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2315_c7_37fa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;

     -- t16_MUX[uxn_opcodes_h_l2315_c7_37fa] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2315_c7_37fa_cond <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_cond;
     t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue;
     t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output := t16_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2312_c7_d7c4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2320_c7_ca68] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output := result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2320_c7_ca68_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2312_c7_d7c4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2315_c7_37fa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2312_c7_d7c4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2315_c7_37fa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;

     -- t16_MUX[uxn_opcodes_h_l2312_c7_d7c4] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond;
     t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue;
     t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output := t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2315_c7_37fa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output := result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2307_c2_96b3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2315_c7_37fa_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2312_c7_d7c4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output := result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2307_c2_96b3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2307_c2_96b3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2312_c7_d7c4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2312_c7_d7c4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;

     -- t16_MUX[uxn_opcodes_h_l2307_c2_96b3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2307_c2_96b3_cond <= VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_cond;
     t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue;
     t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output := t16_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2312_c7_d7c4_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2307_c2_96b3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2307_c2_96b3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2307_c2_96b3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2341_l2303_DUPLICATE_bafb LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2341_l2303_DUPLICATE_bafb_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_25e8(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2307_c2_96b3_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2341_l2303_DUPLICATE_bafb_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l2341_l2303_DUPLICATE_bafb_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
