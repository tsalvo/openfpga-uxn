-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity mul_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_64d180f1;
architecture arch of mul_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1970_c6_8ded]
signal BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal n8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal t8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1970_c2_31ad]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1983_c11_faf6]
signal BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1983_c7_edae]
signal n8_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1983_c7_edae]
signal t8_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1983_c7_edae]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1983_c7_edae]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1983_c7_edae]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1983_c7_edae]
signal result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1983_c7_edae]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1986_c11_250f]
signal BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1986_c7_33b5]
signal n8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1986_c7_33b5]
signal t8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1986_c7_33b5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1986_c7_33b5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1986_c7_33b5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1986_c7_33b5]
signal result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1986_c7_33b5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1989_c11_ae72]
signal BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1989_c7_47ff]
signal n8_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1989_c7_47ff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1989_c7_47ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1989_c7_47ff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1989_c7_47ff]
signal result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1989_c7_47ff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1991_c30_b7fc]
signal sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1994_c21_7ea4]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_return_output : unsigned(15 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a6df( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded
BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_left,
BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_right,
BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output);

-- n8_MUX_uxn_opcodes_h_l1970_c2_31ad
n8_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
n8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- t8_MUX_uxn_opcodes_h_l1970_c2_31ad
t8_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
t8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad
result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad
result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad
result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad
result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad
result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad
result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad
result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6
BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_left,
BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_right,
BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output);

-- n8_MUX_uxn_opcodes_h_l1983_c7_edae
n8_MUX_uxn_opcodes_h_l1983_c7_edae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1983_c7_edae_cond,
n8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue,
n8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse,
n8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output);

-- t8_MUX_uxn_opcodes_h_l1983_c7_edae
t8_MUX_uxn_opcodes_h_l1983_c7_edae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1983_c7_edae_cond,
t8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue,
t8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse,
t8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae
result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae
result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_cond,
result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f
BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_left,
BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_right,
BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output);

-- n8_MUX_uxn_opcodes_h_l1986_c7_33b5
n8_MUX_uxn_opcodes_h_l1986_c7_33b5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond,
n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue,
n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse,
n8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output);

-- t8_MUX_uxn_opcodes_h_l1986_c7_33b5
t8_MUX_uxn_opcodes_h_l1986_c7_33b5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond,
t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue,
t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse,
t8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5
result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5
result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5
result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72
BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_left,
BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_right,
BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output);

-- n8_MUX_uxn_opcodes_h_l1989_c7_47ff
n8_MUX_uxn_opcodes_h_l1989_c7_47ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1989_c7_47ff_cond,
n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue,
n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse,
n8_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff
result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff
result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff
result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_cond,
result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff
result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc
sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_ins,
sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_x,
sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_y,
sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4 : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output,
 n8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 t8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output,
 n8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output,
 t8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output,
 n8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output,
 t8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output,
 n8_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output,
 sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1975_c3_df81 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1980_c3_5d72 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1984_c3_046e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1993_c3_bf4b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l1994_c3_fcc5 : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1986_l1970_l1989_l1983_DUPLICATE_bef2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_1ffe_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_f83a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_2f7e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1986_l1989_DUPLICATE_e50b_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1966_l1998_DUPLICATE_4df5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1984_c3_046e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1984_c3_046e;
     VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1993_c3_bf4b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1993_c3_bf4b;
     VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1980_c3_5d72 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1980_c3_5d72;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1975_c3_df81 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1975_c3_df81;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1970_c6_8ded] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_left;
     BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output := BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1986_c11_250f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output := result.is_vram_write;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1994_c21_7ea4] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output := result.is_ram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_1ffe LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_1ffe_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_f83a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_f83a_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_2f7e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_2f7e_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1986_l1989_DUPLICATE_e50b LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1986_l1989_DUPLICATE_e50b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1983_c11_faf6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1989_c11_ae72] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_left;
     BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output := BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1991_c30_b7fc] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_ins;
     sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_x;
     sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_return_output := sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1986_l1970_l1989_l1983_DUPLICATE_bef2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1986_l1970_l1989_l1983_DUPLICATE_bef2_return_output := result.u8_value;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1970_c6_8ded_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1983_c11_faf6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1986_c11_250f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1989_c11_ae72_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l1994_c3_fcc5 := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1994_c21_7ea4_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_1ffe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_1ffe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_1ffe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_f83a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_f83a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_f83a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_2f7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_2f7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1986_l1989_l1983_DUPLICATE_2f7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1986_l1989_DUPLICATE_e50b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1986_l1989_DUPLICATE_e50b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1986_l1970_l1989_l1983_DUPLICATE_bef2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1986_l1970_l1989_l1983_DUPLICATE_bef2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1986_l1970_l1989_l1983_DUPLICATE_bef2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1986_l1970_l1989_l1983_DUPLICATE_bef2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1970_c2_31ad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1991_c30_b7fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue := VAR_result_u8_value_uxn_opcodes_h_l1994_c3_fcc5;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- t8_MUX[uxn_opcodes_h_l1986_c7_33b5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond;
     t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue;
     t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output := t8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1989_c7_47ff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1989_c7_47ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;

     -- n8_MUX[uxn_opcodes_h_l1989_c7_47ff] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1989_c7_47ff_cond <= VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_cond;
     n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue;
     n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output := n8_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1989_c7_47ff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1989_c7_47ff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output := result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1989_c7_47ff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1989_c7_47ff_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;
     -- t8_MUX[uxn_opcodes_h_l1983_c7_edae] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1983_c7_edae_cond <= VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_cond;
     t8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue;
     t8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output := t8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1986_c7_33b5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1986_c7_33b5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_cond;
     n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue;
     n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output := n8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1986_c7_33b5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1986_c7_33b5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1986_c7_33b5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1986_c7_33b5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1986_c7_33b5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;
     -- n8_MUX[uxn_opcodes_h_l1983_c7_edae] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1983_c7_edae_cond <= VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_cond;
     n8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue;
     n8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output := n8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1983_c7_edae] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_return_output := result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;

     -- t8_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := t8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1983_c7_edae] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1983_c7_edae] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1983_c7_edae] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1983_c7_edae] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1983_c7_edae_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- n8_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := n8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1970_c2_31ad] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output := result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1966_l1998_DUPLICATE_4df5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1966_l1998_DUPLICATE_4df5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a6df(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1970_c2_31ad_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1966_l1998_DUPLICATE_4df5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1966_l1998_DUPLICATE_4df5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
