-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sth2_0CLK_55b6500a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth2_0CLK_55b6500a;
architecture arch of sth2_0CLK_55b6500a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2419_c6_096b]
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2419_c2_36c0]
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_9136]
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2432_c7_95c7]
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2432_c7_95c7]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_95c7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_95c7]
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_95c7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_95c7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_95c7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(3 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2432_c7_95c7]
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_3c5c]
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2435_c7_8f4c]
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2435_c7_8f4c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_8f4c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_8f4c]
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_8f4c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_8f4c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_8f4c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(3 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2435_c7_8f4c]
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2437_c30_9946]
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_ee29]
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2439_c7_2a1b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2439_c7_2a1b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2439_c7_2a1b]
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_2a1b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_2a1b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2439_c7_2a1b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(3 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2439_c7_2a1b]
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2447_c11_8551]
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2447_c7_d2e5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2447_c7_d2e5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2447_c7_d2e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2447_c7_d2e5]
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_ee25( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_left,
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_right,
BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0
t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0
t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_cond,
t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue,
t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse,
t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_left,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_right,
BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7
t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_cond,
t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue,
t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse,
t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7
t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_cond,
t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue,
t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse,
t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_left,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_right,
BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c
t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond,
t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue,
t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse,
t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c
t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond,
t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue,
t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse,
t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2437_c30_9946
sp_relative_shift_uxn_opcodes_h_l2437_c30_9946 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_ins,
sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_x,
sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_y,
sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_left,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_right,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b
t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond,
t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue,
t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse,
t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_left,
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_right,
BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output,
 t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output,
 t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output,
 t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output,
 t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output,
 t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output,
 t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_3a01 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_1950 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_17da : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_dbc3 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_e750 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_2dc8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_10cd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_6b6c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_54e1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_82d7_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_5f0e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_cafe_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_a87c_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2454_l2415_DUPLICATE_a58f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_right := to_unsigned(2, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_e750 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2444_c3_e750;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_3a01 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2424_c3_3a01;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_1950 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2429_c3_1950;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_dbc3 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2442_c3_dbc3;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_10cd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2449_c3_10cd;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_2dc8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2448_c3_2dc8;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_17da := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2433_c3_17da;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_left := VAR_phase;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse := t16_low;
     -- BIN_OP_EQ[uxn_opcodes_h_l2432_c11_9136] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_left;
     BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output := BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2419_c6_096b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_6b6c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_6b6c_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_82d7 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_82d7_return_output := result.sp_relative_shift;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_cafe LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_cafe_return_output := result.is_opc_done;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_ee29] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_left;
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output := BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2447_c11_8551] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_left;
     BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output := BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_54e1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_54e1_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_5f0e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_5f0e_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_a87c LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_a87c_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2435_c11_3c5c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2437_c30_9946] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_ins;
     sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_x;
     sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_return_output := sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c6_096b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2432_c11_9136_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2435_c11_3c5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_ee29_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2447_c11_8551_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_82d7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2432_l2447_DUPLICATE_82d7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_cafe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_cafe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_cafe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2439_l2432_l2447_l2435_DUPLICATE_cafe_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_54e1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_54e1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_54e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_5f0e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_5f0e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2439_l2432_l2435_DUPLICATE_5f0e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_a87c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2447_l2435_DUPLICATE_a87c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_6b6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_6b6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_6b6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2432_l2447_l2435_l2419_DUPLICATE_6b6c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2419_c2_36c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2437_c30_9946_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2447_c7_d2e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_2a1b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2439_c7_2a1b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2447_c7_d2e5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2439_c7_2a1b] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond;
     t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output := t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2447_c7_d2e5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2447_c7_d2e5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2435_c7_8f4c] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond;
     t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output := t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2447_c7_d2e5_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2435_c7_8f4c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2439_c7_2a1b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2439_c7_2a1b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_2a1b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2432_c7_95c7] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_cond;
     t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output := t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2439_c7_2a1b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2435_c7_8f4c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2435_c7_8f4c] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond;
     t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output := t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2439_c7_2a1b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2435_c7_8f4c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2435_c7_8f4c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2435_c7_8f4c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2432_c7_95c7] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_cond;
     t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output := t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2435_c7_8f4c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2432_c7_95c7] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2432_c7_95c7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2435_c7_8f4c_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2432_c7_95c7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2432_c7_95c7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2432_c7_95c7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2432_c7_95c7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2432_c7_95c7_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2419_c2_36c0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2454_l2415_DUPLICATE_a58f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2454_l2415_DUPLICATE_a58f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_ee25(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2419_c2_36c0_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2454_l2415_DUPLICATE_a58f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l2454_l2415_DUPLICATE_a58f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
