-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity neq_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_226c8821;
architecture arch of neq_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1242_c6_7108]
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal n8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1242_c2_e48b]
signal t8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1255_c11_438b]
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1255_c7_d8a0]
signal n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1255_c7_d8a0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1255_c7_d8a0]
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1255_c7_d8a0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1255_c7_d8a0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1255_c7_d8a0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1255_c7_d8a0]
signal t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1258_c11_245f]
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1258_c7_0d6f]
signal n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1258_c7_0d6f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1258_c7_0d6f]
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1258_c7_0d6f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1258_c7_0d6f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1258_c7_0d6f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1258_c7_0d6f]
signal t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1261_c11_80ed]
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1261_c7_ca8b]
signal n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1261_c7_ca8b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1261_c7_ca8b]
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1261_c7_ca8b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1261_c7_ca8b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1261_c7_ca8b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1263_c30_9fe8]
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1266_c21_befa]
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1266_c21_0506]
signal MUX_uxn_opcodes_h_l1266_c21_0506_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_0506_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_0506_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1266_c21_0506_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_left,
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_right,
BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output);

-- n8_MUX_uxn_opcodes_h_l1242_c2_e48b
n8_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
n8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- t8_MUX_uxn_opcodes_h_l1242_c2_e48b
t8_MUX_uxn_opcodes_h_l1242_c2_e48b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond,
t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue,
t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse,
t8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_left,
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_right,
BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output);

-- n8_MUX_uxn_opcodes_h_l1255_c7_d8a0
n8_MUX_uxn_opcodes_h_l1255_c7_d8a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond,
n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue,
n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse,
n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output);

-- t8_MUX_uxn_opcodes_h_l1255_c7_d8a0
t8_MUX_uxn_opcodes_h_l1255_c7_d8a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond,
t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue,
t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse,
t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_left,
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_right,
BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output);

-- n8_MUX_uxn_opcodes_h_l1258_c7_0d6f
n8_MUX_uxn_opcodes_h_l1258_c7_0d6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond,
n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue,
n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse,
n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output);

-- t8_MUX_uxn_opcodes_h_l1258_c7_0d6f
t8_MUX_uxn_opcodes_h_l1258_c7_0d6f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond,
t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue,
t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse,
t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_left,
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_right,
BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output);

-- n8_MUX_uxn_opcodes_h_l1261_c7_ca8b
n8_MUX_uxn_opcodes_h_l1261_c7_ca8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond,
n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue,
n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse,
n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8
sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_ins,
sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_x,
sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_y,
sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_left,
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_right,
BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_return_output);

-- MUX_uxn_opcodes_h_l1266_c21_0506
MUX_uxn_opcodes_h_l1266_c21_0506 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1266_c21_0506_cond,
MUX_uxn_opcodes_h_l1266_c21_0506_iftrue,
MUX_uxn_opcodes_h_l1266_c21_0506_iffalse,
MUX_uxn_opcodes_h_l1266_c21_0506_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output,
 n8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 t8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output,
 n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output,
 t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output,
 n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output,
 t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output,
 n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_return_output,
 MUX_uxn_opcodes_h_l1266_c21_0506_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_50a5 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_ecc5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_0dbe : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_b531 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_0506_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_0506_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_0506_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1266_c21_0506_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_7d98_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_3343_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_72fb_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_2cf1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_e373_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1270_l1238_DUPLICATE_f06a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_ecc5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1252_c3_ecc5;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_0dbe := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1256_c3_0dbe;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_b531 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1265_c3_b531;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_y := resize(to_signed(-1, 2), 4);
     VAR_MUX_uxn_opcodes_h_l1266_c21_0506_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_MUX_uxn_opcodes_h_l1266_c21_0506_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_50a5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1247_c3_50a5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1242_c6_7108] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_left;
     BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output := BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1266_c21_befa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_left;
     BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_return_output := BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1258_c11_245f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l1263_c30_9fe8] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_ins;
     sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_x;
     sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_return_output := sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_7d98 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_7d98_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_72fb LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_72fb_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1255_c11_438b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1261_c11_80ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_3343 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_3343_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_e373 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_e373_return_output := result.stack_address_sp_offset;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_2cf1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_2cf1_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1242_c6_7108_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1255_c11_438b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1258_c11_245f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1261_c11_80ed_return_output;
     VAR_MUX_uxn_opcodes_h_l1266_c21_0506_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1266_c21_befa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_72fb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_72fb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_72fb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_2cf1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_2cf1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_2cf1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_3343_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_3343_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1255_l1258_l1261_DUPLICATE_3343_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_e373_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1258_l1261_DUPLICATE_e373_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_7d98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_7d98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_7d98_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1255_l1258_l1242_l1261_DUPLICATE_7d98_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1242_c2_e48b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1263_c30_9fe8_return_output;
     -- n8_MUX[uxn_opcodes_h_l1261_c7_ca8b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond;
     n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue;
     n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output := n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1258_c7_0d6f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond;
     t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue;
     t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output := t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1261_c7_ca8b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1261_c7_ca8b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1261_c7_ca8b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1261_c7_ca8b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;

     -- MUX[uxn_opcodes_h_l1266_c21_0506] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1266_c21_0506_cond <= VAR_MUX_uxn_opcodes_h_l1266_c21_0506_cond;
     MUX_uxn_opcodes_h_l1266_c21_0506_iftrue <= VAR_MUX_uxn_opcodes_h_l1266_c21_0506_iftrue;
     MUX_uxn_opcodes_h_l1266_c21_0506_iffalse <= VAR_MUX_uxn_opcodes_h_l1266_c21_0506_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1266_c21_0506_return_output := MUX_uxn_opcodes_h_l1266_c21_0506_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue := VAR_MUX_uxn_opcodes_h_l1266_c21_0506_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;
     -- t8_MUX[uxn_opcodes_h_l1255_c7_d8a0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond;
     t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue;
     t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output := t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1258_c7_0d6f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1258_c7_0d6f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond;
     n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue;
     n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output := n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1258_c7_0d6f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1258_c7_0d6f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1261_c7_ca8b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1258_c7_0d6f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1261_c7_ca8b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;
     -- t8_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := t8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1255_c7_d8a0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1258_c7_0d6f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1255_c7_d8a0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1255_c7_d8a0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;

     -- n8_MUX[uxn_opcodes_h_l1255_c7_d8a0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond;
     n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue;
     n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output := n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1255_c7_d8a0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1258_c7_0d6f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1255_c7_d8a0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;

     -- n8_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := n8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1255_c7_d8a0_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1242_c2_e48b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1270_l1238_DUPLICATE_f06a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1270_l1238_DUPLICATE_f06a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1242_c2_e48b_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1270_l1238_DUPLICATE_f06a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1270_l1238_DUPLICATE_f06a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
