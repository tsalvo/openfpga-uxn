-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity ldz_0CLK_b128164d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_b128164d;
architecture arch of ldz_0CLK_b128164d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_12da]
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(15 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1437_c2_8f5f]
signal t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_0291]
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1450_c7_609f]
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_609f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1450_c7_609f]
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_609f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1450_c7_609f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1450_c7_609f]
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_609f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1450_c7_609f]
signal t8_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1453_c11_5a35]
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1453_c7_109a]
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1453_c7_109a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1453_c7_109a]
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1453_c7_109a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1453_c7_109a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1453_c7_109a]
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1453_c7_109a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1453_c7_109a]
signal t8_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1455_c30_a36e]
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1458_c11_998f]
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1458_c7_e6da]
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1458_c7_e6da]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1458_c7_e6da]
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1458_c7_e6da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1458_c7_e6da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1458_c7_e6da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1461_c11_1854]
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1461_c7_49a4]
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1461_c7_49a4]
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1461_c7_49a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1461_c7_49a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1461_c7_49a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_6145( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.u16_value := ref_toks_6;
      base.is_stack_index_flipped := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_opc_done := ref_toks_9;
      base.stack_address_sp_offset := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_left,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_right,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f
tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- t8_MUX_uxn_opcodes_h_l1437_c2_8f5f
t8_MUX_uxn_opcodes_h_l1437_c2_8f5f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond,
t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue,
t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse,
t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_left,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_right,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1450_c7_609f
tmp8_MUX_uxn_opcodes_h_l1450_c7_609f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_cond,
tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue,
tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse,
tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_return_output);

-- t8_MUX_uxn_opcodes_h_l1450_c7_609f
t8_MUX_uxn_opcodes_h_l1450_c7_609f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1450_c7_609f_cond,
t8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue,
t8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse,
t8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_left,
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_right,
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1453_c7_109a
tmp8_MUX_uxn_opcodes_h_l1453_c7_109a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_cond,
tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue,
tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse,
tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_return_output);

-- t8_MUX_uxn_opcodes_h_l1453_c7_109a
t8_MUX_uxn_opcodes_h_l1453_c7_109a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1453_c7_109a_cond,
t8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue,
t8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse,
t8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e
sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_ins,
sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_x,
sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_y,
sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_left,
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_right,
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da
tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_cond,
tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue,
tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse,
tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_cond,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_left,
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_right,
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4
tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_cond,
tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue,
tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse,
tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output,
 tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output,
 tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_return_output,
 t8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output,
 tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_return_output,
 t8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output,
 sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output,
 tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output,
 tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_8622 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_2c4a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_7415 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_88c9_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_053c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_29b4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1458_l1453_l1450_l1437_l1461_DUPLICATE_6c9c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_744b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_b290_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_cc74_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_4e15_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_9f59_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l1469_l1433_DUPLICATE_90a8_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_8622 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_8622;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_right := to_unsigned(2, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_2c4a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_2c4a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_7415 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_7415;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_053c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_053c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_29b4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_29b4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_right := to_unsigned(4, 3);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse := tmp8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_b290 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_b290_return_output := result.is_opc_done;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1456_c22_88c9] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_88c9_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1455_c30_a36e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_ins;
     sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_x;
     sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_return_output := sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1461_c11_1854] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_left;
     BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output := BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1453_c11_5a35] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_left;
     BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output := BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_12da] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_left;
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output := BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1458_c11_998f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output := result.is_ram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_4e15 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_4e15_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_0291] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_left;
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output := BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_744b LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_744b_return_output := result.u16_value;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1458_l1453_l1450_l1437_l1461_DUPLICATE_6c9c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1458_l1453_l1450_l1437_l1461_DUPLICATE_6c9c_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_9f59 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_9f59_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_cc74 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_cc74_return_output := result.is_stack_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_12da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0291_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_5a35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_998f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_1854_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_88c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_4e15_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_4e15_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_744b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_744b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_744b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_b290_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_b290_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_b290_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_b290_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_cc74_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_cc74_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_cc74_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_cc74_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_9f59_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_9f59_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_9f59_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1458_l1453_l1450_l1437_l1461_DUPLICATE_6c9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1458_l1453_l1450_l1437_l1461_DUPLICATE_6c9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1458_l1453_l1450_l1437_l1461_DUPLICATE_6c9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1458_l1453_l1450_l1437_l1461_DUPLICATE_6c9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1458_l1453_l1450_l1437_l1461_DUPLICATE_6c9c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_8f5f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_a36e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1461_c7_49a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1461_c7_49a4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1458_c7_e6da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1453_c7_109a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output := result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1461_c7_49a4] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_cond;
     tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output := tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1461_c7_49a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1453_c7_109a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1453_c7_109a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_cond;
     t8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue;
     t8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output := t8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1461_c7_49a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_49a4_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1458_c7_e6da] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_cond;
     tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output := tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;

     -- t8_MUX[uxn_opcodes_h_l1450_c7_609f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1450_c7_609f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_cond;
     t8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue;
     t8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output := t8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1458_c7_e6da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1458_c7_e6da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1450_c7_609f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output := result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1453_c7_109a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1458_c7_e6da] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output := result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1458_c7_e6da] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_e6da_return_output;
     -- t8_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1453_c7_109a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1453_c7_109a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1453_c7_109a] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_cond;
     tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output := tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1453_c7_109a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1450_c7_609f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1453_c7_109a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_109a_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_609f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1450_c7_609f] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_cond;
     tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output := tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1450_c7_609f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_609f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_609f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_609f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_8f5f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l1469_l1433_DUPLICATE_90a8 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l1469_l1433_DUPLICATE_90a8_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_6145(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_8f5f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l1469_l1433_DUPLICATE_90a8_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_6145_uxn_opcodes_h_l1469_l1433_DUPLICATE_90a8_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
