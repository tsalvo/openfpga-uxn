-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity lth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_226c8821;
architecture arch of lth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1912_c6_935d]
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal n8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal t8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1912_c2_efe6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1925_c11_ea3f]
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1925_c7_5992]
signal n8_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1925_c7_5992]
signal t8_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1925_c7_5992]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1925_c7_5992]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1925_c7_5992]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1925_c7_5992]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1925_c7_5992]
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1928_c11_d940]
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1928_c7_6891]
signal n8_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1928_c7_6891]
signal t8_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1928_c7_6891]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1928_c7_6891]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1928_c7_6891]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1928_c7_6891]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1928_c7_6891]
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1931_c11_e648]
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1931_c7_c362]
signal n8_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1931_c7_c362]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1931_c7_c362]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1931_c7_c362]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1931_c7_c362]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1931_c7_c362]
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1933_c30_561e]
signal sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1936_c21_4800]
signal BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1936_c21_8a13]
signal MUX_uxn_opcodes_h_l1936_c21_8a13_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1936_c21_8a13_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1936_c21_8a13_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1936_c21_8a13_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e848( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d
BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_left,
BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_right,
BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output);

-- n8_MUX_uxn_opcodes_h_l1912_c2_efe6
n8_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
n8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- t8_MUX_uxn_opcodes_h_l1912_c2_efe6
t8_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
t8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_left,
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_right,
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output);

-- n8_MUX_uxn_opcodes_h_l1925_c7_5992
n8_MUX_uxn_opcodes_h_l1925_c7_5992 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1925_c7_5992_cond,
n8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue,
n8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse,
n8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output);

-- t8_MUX_uxn_opcodes_h_l1925_c7_5992
t8_MUX_uxn_opcodes_h_l1925_c7_5992 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1925_c7_5992_cond,
t8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue,
t8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse,
t8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_cond,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_left,
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_right,
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output);

-- n8_MUX_uxn_opcodes_h_l1928_c7_6891
n8_MUX_uxn_opcodes_h_l1928_c7_6891 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1928_c7_6891_cond,
n8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue,
n8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse,
n8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output);

-- t8_MUX_uxn_opcodes_h_l1928_c7_6891
t8_MUX_uxn_opcodes_h_l1928_c7_6891 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1928_c7_6891_cond,
t8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue,
t8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse,
t8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_cond,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_left,
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_right,
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output);

-- n8_MUX_uxn_opcodes_h_l1931_c7_c362
n8_MUX_uxn_opcodes_h_l1931_c7_c362 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1931_c7_c362_cond,
n8_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue,
n8_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse,
n8_MUX_uxn_opcodes_h_l1931_c7_c362_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_cond,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1933_c30_561e
sp_relative_shift_uxn_opcodes_h_l1933_c30_561e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_ins,
sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_x,
sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_y,
sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800
BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_left,
BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_right,
BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_return_output);

-- MUX_uxn_opcodes_h_l1936_c21_8a13
MUX_uxn_opcodes_h_l1936_c21_8a13 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1936_c21_8a13_cond,
MUX_uxn_opcodes_h_l1936_c21_8a13_iftrue,
MUX_uxn_opcodes_h_l1936_c21_8a13_iffalse,
MUX_uxn_opcodes_h_l1936_c21_8a13_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output,
 n8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 t8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output,
 n8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output,
 t8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output,
 n8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output,
 t8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output,
 n8_MUX_uxn_opcodes_h_l1931_c7_c362_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_return_output,
 sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_return_output,
 MUX_uxn_opcodes_h_l1936_c21_8a13_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1917_c3_c4fc : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_58f9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_f5e2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1935_c3_4f49 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1912_l1928_l1931_DUPLICATE_3c69_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_f17c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_41da_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_19a7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1928_l1931_DUPLICATE_9b41_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1940_l1908_DUPLICATE_6edf_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_f5e2 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_f5e2;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_58f9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_58f9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1935_c3_4f49 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1935_c3_4f49;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1917_c3_c4fc := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1917_c3_c4fc;
     VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_right := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_y := resize(to_signed(-1, 2), 4);
     VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1925_c11_ea3f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output := result.is_stack_index_flipped;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1928_l1931_DUPLICATE_9b41 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1928_l1931_DUPLICATE_9b41_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1928_c11_d940] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_left;
     BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output := BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_41da LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_41da_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1912_c6_935d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;

     -- BIN_OP_LT[uxn_opcodes_h_l1936_c21_4800] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_left;
     BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_return_output := BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1912_l1928_l1931_DUPLICATE_3c69 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1912_l1928_l1931_DUPLICATE_3c69_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_f17c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_f17c_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1933_c30_561e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_ins;
     sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_x;
     sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_return_output := sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output := result.is_ram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1931_c11_e648] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_left;
     BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output := BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_19a7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_19a7_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_935d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ea3f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_d940_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_e648_return_output;
     VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_4800_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_41da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_41da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_41da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_19a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_19a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_19a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_f17c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_f17c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1928_l1931_DUPLICATE_f17c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1928_l1931_DUPLICATE_9b41_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1928_l1931_DUPLICATE_9b41_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1912_l1928_l1931_DUPLICATE_3c69_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1912_l1928_l1931_DUPLICATE_3c69_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1912_l1928_l1931_DUPLICATE_3c69_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1912_l1928_l1931_DUPLICATE_3c69_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1912_c2_efe6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_561e_return_output;
     -- t8_MUX[uxn_opcodes_h_l1928_c7_6891] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1928_c7_6891_cond <= VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_cond;
     t8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue;
     t8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output := t8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1931_c7_c362] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1931_c7_c362] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- n8_MUX[uxn_opcodes_h_l1931_c7_c362] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1931_c7_c362_cond <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_cond;
     n8_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue;
     n8_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_return_output := n8_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;

     -- MUX[uxn_opcodes_h_l1936_c21_8a13] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1936_c21_8a13_cond <= VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_cond;
     MUX_uxn_opcodes_h_l1936_c21_8a13_iftrue <= VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_iftrue;
     MUX_uxn_opcodes_h_l1936_c21_8a13_iffalse <= VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_return_output := MUX_uxn_opcodes_h_l1936_c21_8a13_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1931_c7_c362] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1931_c7_c362] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue := VAR_MUX_uxn_opcodes_h_l1936_c21_8a13_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;
     -- t8_MUX[uxn_opcodes_h_l1925_c7_5992] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1925_c7_5992_cond <= VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_cond;
     t8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue;
     t8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output := t8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1928_c7_6891] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1928_c7_6891] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1931_c7_c362] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_return_output := result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;

     -- n8_MUX[uxn_opcodes_h_l1928_c7_6891] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1928_c7_6891_cond <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_cond;
     n8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue;
     n8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output := n8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1928_c7_6891] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1928_c7_6891] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_c362_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1925_c7_5992] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;

     -- n8_MUX[uxn_opcodes_h_l1925_c7_5992] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1925_c7_5992_cond <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_cond;
     n8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue;
     n8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output := n8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1925_c7_5992] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1928_c7_6891] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_return_output := result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1925_c7_5992] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;

     -- t8_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := t8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1925_c7_5992] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_6891_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;
     -- n8_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := n8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1925_c7_5992] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_return_output := result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5992_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1912_c2_efe6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1940_l1908_DUPLICATE_6edf LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1940_l1908_DUPLICATE_6edf_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e848(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_efe6_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1940_l1908_DUPLICATE_6edf_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1940_l1908_DUPLICATE_6edf_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
