-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity stz2_0CLK_75b4bee3 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end stz2_0CLK_75b4bee3;
architecture arch of stz2_0CLK_75b4bee3 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n16_low : unsigned(7 downto 0);
signal REG_COMB_n16_high : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1557_c6_8c8c]
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l1557_c2_2566]
signal n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1557_c2_2566]
signal t8_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1557_c2_2566]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1557_c2_2566]
signal n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1570_c11_a830]
signal BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1570_c7_2f2e]
signal n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1573_c11_e01c]
signal BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal t8_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1573_c7_cb91]
signal n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1577_c11_522a]
signal BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l1577_c7_f035]
signal n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1577_c7_f035]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1577_c7_f035]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1577_c7_f035]
signal result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1577_c7_f035]
signal result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1577_c7_f035]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(0 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1577_c7_f035]
signal n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1579_c30_1227]
signal sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1584_c11_de1b]
signal BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1584_c7_0a47]
signal result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1584_c7_0a47]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1584_c7_0a47]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1584_c7_0a47]
signal result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : unsigned(7 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l1584_c7_0a47]
signal n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1587_c33_e8b4]
signal BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_return_output : unsigned(8 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint9_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(8 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_1899( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_index_flipped := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.u16_value := ref_toks_8;
      base.is_ram_write := ref_toks_9;
      base.stack_address_sp_offset := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_left,
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_right,
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output);

-- n16_high_MUX_uxn_opcodes_h_l1557_c2_2566
n16_high_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- t8_MUX_uxn_opcodes_h_l1557_c2_2566
t8_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
t8_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
t8_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
t8_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566
result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566
result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566
result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566
result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566
result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1557_c2_2566
n16_low_MUX_uxn_opcodes_h_l1557_c2_2566 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_cond,
n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue,
n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse,
n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830
BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_left,
BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_right,
BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output);

-- n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e
n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- t8_MUX_uxn_opcodes_h_l1570_c7_2f2e
t8_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e
result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e
result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e
result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e
result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e
n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond,
n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue,
n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse,
n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c
BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_left,
BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_right,
BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output);

-- n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91
n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- t8_MUX_uxn_opcodes_h_l1573_c7_cb91
t8_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
t8_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91
result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91
result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91
result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91
result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91
result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91
n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_cond,
n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue,
n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse,
n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a
BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_left,
BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_right,
BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output);

-- n16_high_MUX_uxn_opcodes_h_l1577_c7_f035
n16_high_MUX_uxn_opcodes_h_l1577_c7_f035 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_cond,
n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue,
n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse,
n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035
result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035
result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond,
result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035
result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond,
result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035
result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1577_c7_f035
n16_low_MUX_uxn_opcodes_h_l1577_c7_f035 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_cond,
n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue,
n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse,
n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1579_c30_1227
sp_relative_shift_uxn_opcodes_h_l1579_c30_1227 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_ins,
sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_x,
sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_y,
sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b
BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_left,
BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_right,
BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47
result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond,
result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47
result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47
result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47
result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond,
result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output);

-- n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47
n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_cond,
n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue,
n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse,
n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4
BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_left,
BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_right,
BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n16_low,
 n16_high,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output,
 n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 t8_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output,
 n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output,
 n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 t8_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output,
 n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_return_output,
 n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_return_output,
 sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output,
 n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1562_c3_5f98 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1567_c3_c998 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1571_c3_e0d3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1575_c3_5d38 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1573_c7_cb91_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1581_c22_f3ee_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1586_c3_b1ef : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_return_output : unsigned(8 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1587_c22_6378_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_c895_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_21ef_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1570_l1573_l1584_DUPLICATE_e53d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1570_l1577_l1573_l1584_DUPLICATE_8d33_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1570_l1577_l1573_DUPLICATE_2457_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1899_uxn_opcodes_h_l1592_l1552_DUPLICATE_025f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n16_low : unsigned(7 downto 0);
variable REG_VAR_n16_high : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n16_low := n16_low;
  REG_VAR_n16_high := n16_high;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_y := resize(to_signed(-3, 3), 4);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1562_c3_5f98 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1562_c3_5f98;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_right := to_unsigned(4, 3);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1567_c3_c998 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1567_c3_c998;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1586_c3_b1ef := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1586_c3_b1ef;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1575_c3_5d38 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1575_c3_5d38;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1571_c3_e0d3 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1571_c3_e0d3;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_ins := VAR_ins;
     VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse := n16_high;
     VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse := n16_low;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_left := VAR_phase;
     VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue := VAR_previous_stack_read;
     VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := t8;
     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_21ef LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_21ef_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1584_c11_de1b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1557_c2_2566_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1570_l1577_l1573_DUPLICATE_2457 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1570_l1577_l1573_DUPLICATE_2457_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1577_c11_522a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_c895 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_c895_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l1579_c30_1227] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_ins;
     sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_x;
     sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_return_output := sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1570_l1577_l1573_l1584_DUPLICATE_8d33 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1570_l1577_l1573_l1584_DUPLICATE_8d33_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1573_c7_cb91_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1557_c6_8c8c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1557_c2_2566_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1557_c2_2566_return_output := result.is_vram_write;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1587_c33_e8b4] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1573_c11_e01c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1570_l1573_l1584_DUPLICATE_e53d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1570_l1573_l1584_DUPLICATE_e53d_return_output := result.sp_relative_shift;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1581_c22_f3ee] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1581_c22_f3ee_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1557_c2_2566_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1570_c11_a830] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_left;
     BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output := BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;

     -- Submodule level 1
     VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_8c8c_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1570_c11_a830_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1573_c11_e01c_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1577_c11_522a_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1584_c11_de1b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1581_c22_f3ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1570_l1573_l1584_DUPLICATE_e53d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1570_l1573_l1584_DUPLICATE_e53d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1570_l1573_l1584_DUPLICATE_e53d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_21ef_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_21ef_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_21ef_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_21ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1570_l1577_l1573_l1584_DUPLICATE_8d33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1570_l1577_l1573_l1584_DUPLICATE_8d33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1570_l1577_l1573_l1584_DUPLICATE_8d33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1570_l1577_l1573_l1584_DUPLICATE_8d33_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1570_l1577_l1573_DUPLICATE_2457_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1570_l1577_l1573_DUPLICATE_2457_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1570_l1577_l1573_DUPLICATE_2457_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_c895_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_c895_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_c895_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1570_l1573_l1557_l1584_DUPLICATE_c895_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1557_c2_2566_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1557_c2_2566_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1557_c2_2566_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1557_c2_2566_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1573_c7_cb91_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1579_c30_1227_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1577_c7_f035] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- t8_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := t8_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1584_c7_0a47] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output := result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1584_c7_0a47] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l1577_c7_f035] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_cond;
     n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue;
     n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_return_output := n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1584_c7_0a47] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l1584_c7_0a47] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_cond;
     n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output := n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1587_c22_6378] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1587_c22_6378_return_output := CAST_TO_uint16_t_uint9_t(
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1587_c33_e8b4_return_output);

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1587_c22_6378_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- t8_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1584_c7_0a47] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output := result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1577_c7_f035] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l1577_c7_f035] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_cond;
     n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_return_output := n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1577_c7_f035] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output := result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1577_c7_f035] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;

     -- Submodule level 3
     VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1584_c7_0a47_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     -- n16_high_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1577_c7_f035] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output := result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- t8_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     t8_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     t8_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := t8_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- Submodule level 4
     VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1577_c7_f035_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1573_c7_cb91] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output := result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- Submodule level 5
     REG_VAR_n16_high := VAR_n16_high_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1573_c7_cb91_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     -- n16_low_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1570_c7_2f2e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output := result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- Submodule level 6
     REG_VAR_n16_low := VAR_n16_low_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1570_c7_2f2e_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l1557_c2_2566] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output := result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_1899_uxn_opcodes_h_l1592_l1552_DUPLICATE_025f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1899_uxn_opcodes_h_l1592_l1552_DUPLICATE_025f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_1899(
     result,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1557_c2_2566_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_2566_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1899_uxn_opcodes_h_l1592_l1552_DUPLICATE_025f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1899_uxn_opcodes_h_l1592_l1552_DUPLICATE_025f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n16_low <= REG_VAR_n16_low;
REG_COMB_n16_high <= REG_VAR_n16_high;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n16_low <= REG_COMB_n16_low;
     n16_high <= REG_COMB_n16_high;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
