-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity mul_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_bacf6a1d;
architecture arch of mul_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1874_c6_2ed4]
signal BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1874_c1_330d]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1874_c2_f260]
signal n8_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1874_c2_f260]
signal t8_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1874_c2_f260]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1874_c2_f260]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1874_c2_f260]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1874_c2_f260]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1874_c2_f260]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1874_c2_f260]
signal result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1875_c3_038c[uxn_opcodes_h_l1875_c3_038c]
signal printf_uxn_opcodes_h_l1875_c3_038c_uxn_opcodes_h_l1875_c3_038c_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1879_c11_394e]
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1879_c7_c735]
signal n8_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1879_c7_c735]
signal t8_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1879_c7_c735]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1879_c7_c735]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1879_c7_c735]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1879_c7_c735]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1879_c7_c735]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1879_c7_c735]
signal result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1882_c11_4e02]
signal BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1882_c7_2ea9]
signal n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1882_c7_2ea9]
signal t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1882_c7_2ea9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1882_c7_2ea9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1882_c7_2ea9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1882_c7_2ea9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1882_c7_2ea9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1882_c7_2ea9]
signal result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1885_c11_3b81]
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1885_c7_fc04]
signal n8_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1885_c7_fc04]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1885_c7_fc04]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1885_c7_fc04]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1885_c7_fc04]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1885_c7_fc04]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1885_c7_fc04]
signal result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1888_c30_1e0e]
signal sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1891_c21_0114]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1893_c11_1cd8]
signal BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1893_c7_c7ee]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1893_c7_c7ee]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1893_c7_c7ee]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4
BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_left,
BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_right,
BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_return_output);

-- n8_MUX_uxn_opcodes_h_l1874_c2_f260
n8_MUX_uxn_opcodes_h_l1874_c2_f260 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1874_c2_f260_cond,
n8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue,
n8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse,
n8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

-- t8_MUX_uxn_opcodes_h_l1874_c2_f260
t8_MUX_uxn_opcodes_h_l1874_c2_f260 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1874_c2_f260_cond,
t8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue,
t8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse,
t8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_cond,
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

-- printf_uxn_opcodes_h_l1875_c3_038c_uxn_opcodes_h_l1875_c3_038c
printf_uxn_opcodes_h_l1875_c3_038c_uxn_opcodes_h_l1875_c3_038c : entity work.printf_uxn_opcodes_h_l1875_c3_038c_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1875_c3_038c_uxn_opcodes_h_l1875_c3_038c_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_left,
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_right,
BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output);

-- n8_MUX_uxn_opcodes_h_l1879_c7_c735
n8_MUX_uxn_opcodes_h_l1879_c7_c735 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1879_c7_c735_cond,
n8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue,
n8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse,
n8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output);

-- t8_MUX_uxn_opcodes_h_l1879_c7_c735
t8_MUX_uxn_opcodes_h_l1879_c7_c735 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1879_c7_c735_cond,
t8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue,
t8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse,
t8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_cond,
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02
BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_left,
BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_right,
BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output);

-- n8_MUX_uxn_opcodes_h_l1882_c7_2ea9
n8_MUX_uxn_opcodes_h_l1882_c7_2ea9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond,
n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue,
n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse,
n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output);

-- t8_MUX_uxn_opcodes_h_l1882_c7_2ea9
t8_MUX_uxn_opcodes_h_l1882_c7_2ea9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond,
t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue,
t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse,
t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_left,
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_right,
BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output);

-- n8_MUX_uxn_opcodes_h_l1885_c7_fc04
n8_MUX_uxn_opcodes_h_l1885_c7_fc04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1885_c7_fc04_cond,
n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue,
n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse,
n8_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_cond,
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e
sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_ins,
sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_x,
sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_y,
sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114 : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8
BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_left,
BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_right,
BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_return_output,
 n8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
 t8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output,
 n8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output,
 t8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output,
 n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output,
 t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output,
 n8_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output,
 sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1876_c3_187b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1875_c3_038c_uxn_opcodes_h_l1875_c3_038c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1880_c3_a4e5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1890_c3_0dd9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l1891_c3_0f56 : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_8a93_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_81e8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1882_l1885_l1879_l1893_DUPLICATE_ae5c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1882_l1885_DUPLICATE_7cb2_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1870_l1899_DUPLICATE_43cf_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1876_c3_187b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1876_c3_187b;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iffalse := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1890_c3_0dd9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1890_c3_0dd9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1880_c3_a4e5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1880_c3_a4e5;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse := t8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b3_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1893_c11_1cd8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_left;
     BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output := BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1891_c21_0114] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_8a93 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_8a93_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1888_c30_1e0e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_ins;
     sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_x;
     sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_return_output := sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1879_c11_394e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1882_l1885_l1879_l1893_DUPLICATE_ae5c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1882_l1885_l1879_l1893_DUPLICATE_ae5c_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1874_c6_2ed4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1885_c11_3b81] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_left;
     BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output := BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1882_c11_4e02] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_left;
     BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output := BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_81e8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_81e8_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1882_l1885_DUPLICATE_7cb2 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1882_l1885_DUPLICATE_7cb2_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b5_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1874_c6_2ed4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1879_c11_394e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1882_c11_4e02_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1885_c11_3b81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1893_c11_1cd8_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l1891_c3_0f56 := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1891_c21_0114_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1882_l1885_l1879_l1893_DUPLICATE_ae5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1882_l1885_l1879_l1893_DUPLICATE_ae5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1882_l1885_l1879_l1893_DUPLICATE_ae5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1882_l1885_l1879_l1893_DUPLICATE_ae5c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_81e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_81e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_81e8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_81e8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_8a93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_8a93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_8a93_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1882_l1874_l1879_l1893_DUPLICATE_8a93_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1882_l1885_DUPLICATE_7cb2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1882_l1885_DUPLICATE_7cb2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1882_l1874_l1885_l1879_DUPLICATE_c8b3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1888_c30_1e0e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue := VAR_result_u8_value_uxn_opcodes_h_l1891_c3_0f56;
     -- t8_MUX[uxn_opcodes_h_l1882_c7_2ea9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond <= VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond;
     t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue;
     t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output := t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1874_c1_330d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1885_c7_fc04] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1893_c7_c7ee] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1885_c7_fc04] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1885_c7_fc04] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output := result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1893_c7_c7ee] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1893_c7_c7ee] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output;

     -- n8_MUX[uxn_opcodes_h_l1885_c7_fc04] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1885_c7_fc04_cond <= VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_cond;
     n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue;
     n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output := n8_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1875_c3_038c_uxn_opcodes_h_l1875_c3_038c_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1874_c1_330d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1893_c7_c7ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;
     -- t8_MUX[uxn_opcodes_h_l1879_c7_c735] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1879_c7_c735_cond <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_cond;
     t8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue;
     t8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output := t8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1882_c7_2ea9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1885_c7_fc04] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1885_c7_fc04] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1882_c7_2ea9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;

     -- n8_MUX[uxn_opcodes_h_l1882_c7_2ea9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond <= VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond;
     n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue;
     n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output := n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1885_c7_fc04] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;

     -- printf_uxn_opcodes_h_l1875_c3_038c[uxn_opcodes_h_l1875_c3_038c] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1875_c3_038c_uxn_opcodes_h_l1875_c3_038c_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1875_c3_038c_uxn_opcodes_h_l1875_c3_038c_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1882_c7_2ea9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1885_c7_fc04_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1879_c7_c735] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_return_output := result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1882_c7_2ea9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1882_c7_2ea9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1874_c2_f260] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1874_c2_f260_cond <= VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_cond;
     t8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue;
     t8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output := t8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1882_c7_2ea9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1879_c7_c735] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;

     -- n8_MUX[uxn_opcodes_h_l1879_c7_c735] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1879_c7_c735_cond <= VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_cond;
     n8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue;
     n8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output := n8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1879_c7_c735] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1882_c7_2ea9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1874_c2_f260] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;

     -- n8_MUX[uxn_opcodes_h_l1874_c2_f260] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1874_c2_f260_cond <= VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_cond;
     n8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue;
     n8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output := n8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1874_c2_f260] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1879_c7_c735] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1874_c2_f260] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_return_output := result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1879_c7_c735] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1879_c7_c735] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1879_c7_c735_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1874_c2_f260] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1874_c2_f260] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1874_c2_f260] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1870_l1899_DUPLICATE_43cf LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1870_l1899_DUPLICATE_43cf_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b93(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1874_c2_f260_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1874_c2_f260_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1870_l1899_DUPLICATE_43cf_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1870_l1899_DUPLICATE_43cf_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
