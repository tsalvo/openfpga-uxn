-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity lth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_226c8821;
architecture arch of lth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1906_c6_8ee9]
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal t8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal n8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1906_c2_ad15]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1919_c11_161b]
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1919_c7_fa78]
signal t8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1919_c7_fa78]
signal n8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1919_c7_fa78]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1919_c7_fa78]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1919_c7_fa78]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1919_c7_fa78]
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1919_c7_fa78]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1922_c11_261a]
signal BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1922_c7_f8e1]
signal t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1922_c7_f8e1]
signal n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1922_c7_f8e1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1922_c7_f8e1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1922_c7_f8e1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1922_c7_f8e1]
signal result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1922_c7_f8e1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1925_c11_d653]
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1925_c7_3362]
signal n8_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1925_c7_3362]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1925_c7_3362]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1925_c7_3362]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1925_c7_3362]
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1925_c7_3362]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1927_c30_45bd]
signal sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1930_c21_3a26]
signal BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1930_c21_a384]
signal MUX_uxn_opcodes_h_l1930_c21_a384_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1930_c21_a384_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1930_c21_a384_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1930_c21_a384_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_188e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_ram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9
BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_left,
BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_right,
BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output);

-- t8_MUX_uxn_opcodes_h_l1906_c2_ad15
t8_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
t8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- n8_MUX_uxn_opcodes_h_l1906_c2_ad15
n8_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
n8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b
BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_left,
BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_right,
BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output);

-- t8_MUX_uxn_opcodes_h_l1919_c7_fa78
t8_MUX_uxn_opcodes_h_l1919_c7_fa78 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond,
t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue,
t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse,
t8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output);

-- n8_MUX_uxn_opcodes_h_l1919_c7_fa78
n8_MUX_uxn_opcodes_h_l1919_c7_fa78 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond,
n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue,
n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse,
n8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_cond,
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a
BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_left,
BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_right,
BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output);

-- t8_MUX_uxn_opcodes_h_l1922_c7_f8e1
t8_MUX_uxn_opcodes_h_l1922_c7_f8e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond,
t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue,
t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse,
t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output);

-- n8_MUX_uxn_opcodes_h_l1922_c7_f8e1
n8_MUX_uxn_opcodes_h_l1922_c7_f8e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond,
n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue,
n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse,
n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_left,
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_right,
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output);

-- n8_MUX_uxn_opcodes_h_l1925_c7_3362
n8_MUX_uxn_opcodes_h_l1925_c7_3362 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1925_c7_3362_cond,
n8_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue,
n8_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse,
n8_MUX_uxn_opcodes_h_l1925_c7_3362_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_cond,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd
sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_ins,
sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_x,
sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_y,
sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26
BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_left,
BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_right,
BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_return_output);

-- MUX_uxn_opcodes_h_l1930_c21_a384
MUX_uxn_opcodes_h_l1930_c21_a384 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1930_c21_a384_cond,
MUX_uxn_opcodes_h_l1930_c21_a384_iftrue,
MUX_uxn_opcodes_h_l1930_c21_a384_iffalse,
MUX_uxn_opcodes_h_l1930_c21_a384_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output,
 t8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 n8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output,
 t8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output,
 n8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output,
 t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output,
 n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output,
 n8_MUX_uxn_opcodes_h_l1925_c7_3362_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_return_output,
 sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_return_output,
 MUX_uxn_opcodes_h_l1930_c21_a384_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1911_c3_10a7 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1916_c3_a5d7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1920_c3_97e9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_3940 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1930_c21_a384_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1930_c21_a384_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1930_c21_a384_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1930_c21_a384_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1919_l1922_l1906_DUPLICATE_5dad_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_1619_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_cd14_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_c788_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_3868_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1934_l1902_DUPLICATE_7088_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1930_c21_a384_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_3940 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_3940;
     VAR_MUX_uxn_opcodes_h_l1930_c21_a384_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1911_c3_10a7 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1911_c3_10a7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1916_c3_a5d7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1916_c3_a5d7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1920_c3_97e9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1920_c3_97e9;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse := t8;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l1927_c30_45bd] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_ins;
     sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_x;
     sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_return_output := sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1925_c11_d653] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_left;
     BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output := BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_1619 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_1619_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1919_l1922_l1906_DUPLICATE_5dad LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1919_l1922_l1906_DUPLICATE_5dad_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_3868 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_3868_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_c788 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_c788_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1919_c11_161b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output;

     -- BIN_OP_LT[uxn_opcodes_h_l1930_c21_3a26] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_left;
     BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_return_output := BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1906_c6_8ee9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1922_c11_261a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_cd14 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_cd14_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output := result.is_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_8ee9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_161b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_261a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_d653_return_output;
     VAR_MUX_uxn_opcodes_h_l1930_c21_a384_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_3a26_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_1619_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_1619_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_1619_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_c788_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_c788_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_c788_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_cd14_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_cd14_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_cd14_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_3868_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_3868_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1919_l1922_l1906_DUPLICATE_5dad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1919_l1922_l1906_DUPLICATE_5dad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1919_l1922_l1906_DUPLICATE_5dad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1925_l1919_l1922_l1906_DUPLICATE_5dad_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1906_c2_ad15_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_45bd_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- n8_MUX[uxn_opcodes_h_l1925_c7_3362] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1925_c7_3362_cond <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_cond;
     n8_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue;
     n8_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_return_output := n8_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1925_c7_3362] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1925_c7_3362] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1925_c7_3362] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1925_c7_3362] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;

     -- t8_MUX[uxn_opcodes_h_l1922_c7_f8e1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond <= VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond;
     t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue;
     t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output := t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- MUX[uxn_opcodes_h_l1930_c21_a384] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1930_c21_a384_cond <= VAR_MUX_uxn_opcodes_h_l1930_c21_a384_cond;
     MUX_uxn_opcodes_h_l1930_c21_a384_iftrue <= VAR_MUX_uxn_opcodes_h_l1930_c21_a384_iftrue;
     MUX_uxn_opcodes_h_l1930_c21_a384_iffalse <= VAR_MUX_uxn_opcodes_h_l1930_c21_a384_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1930_c21_a384_return_output := MUX_uxn_opcodes_h_l1930_c21_a384_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue := VAR_MUX_uxn_opcodes_h_l1930_c21_a384_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1925_c7_3362] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_return_output := result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1922_c7_f8e1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1919_c7_fa78] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond <= VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond;
     t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue;
     t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output := t8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1922_c7_f8e1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1922_c7_f8e1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1922_c7_f8e1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond;
     n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue;
     n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output := n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1922_c7_f8e1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_3362_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;
     -- n8_MUX[uxn_opcodes_h_l1919_c7_fa78] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond <= VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_cond;
     n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue;
     n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output := n8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1919_c7_fa78] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;

     -- t8_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := t8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1922_c7_f8e1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1919_c7_fa78] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1919_c7_fa78] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1919_c7_fa78] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_f8e1_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- n8_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := n8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1919_c7_fa78] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output := result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_fa78_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1906_c2_ad15] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output := result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1934_l1902_DUPLICATE_7088 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1934_l1902_DUPLICATE_7088_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_188e(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_ad15_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1934_l1902_DUPLICATE_7088_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l1934_l1902_DUPLICATE_7088_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
