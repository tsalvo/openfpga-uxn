-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity inc2_0CLK_180c5210 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_180c5210;
architecture arch of inc2_0CLK_180c5210 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1355_c6_1f9a]
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1355_c2_36cc]
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1368_c11_df5f]
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1368_c7_aa69]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1368_c7_aa69]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1368_c7_aa69]
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1368_c7_aa69]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1368_c7_aa69]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1368_c7_aa69]
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1368_c7_aa69]
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1371_c11_b1b1]
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1371_c7_9acb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1371_c7_9acb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1371_c7_9acb]
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1371_c7_9acb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1371_c7_9acb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1371_c7_9acb]
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1371_c7_9acb]
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1372_c13_5bb4]
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_return_output : unsigned(8 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1373_c30_09f9]
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_0fa0]
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_a19e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c7_a19e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_a19e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_a19e]
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1378_c7_a19e]
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1379_c37_bc63]
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1379_c37_8615]
signal MUX_uxn_opcodes_h_l1379_c37_8615_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_8615_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_8615_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_8615_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1379_c14_6259]
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_left,
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_right,
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc
t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc
t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_cond,
t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue,
t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse,
t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_left,
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_right,
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_cond,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69
t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_cond,
t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue,
t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse,
t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69
t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_cond,
t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue,
t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse,
t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_left,
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_right,
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb
t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_cond,
t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue,
t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse,
t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb
t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_cond,
t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue,
t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse,
t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_left,
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_right,
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9
sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_ins,
sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_x,
sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_y,
sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_left,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_right,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e
t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_cond,
t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue,
t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse,
t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_left,
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_right,
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_return_output);

-- MUX_uxn_opcodes_h_l1379_c37_8615
MUX_uxn_opcodes_h_l1379_c37_8615 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1379_c37_8615_cond,
MUX_uxn_opcodes_h_l1379_c37_8615_iftrue,
MUX_uxn_opcodes_h_l1379_c37_8615_iffalse,
MUX_uxn_opcodes_h_l1379_c37_8615_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259 : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_left,
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_right,
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output,
 t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output,
 t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output,
 t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output,
 t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_return_output,
 sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output,
 t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_return_output,
 MUX_uxn_opcodes_h_l1379_c37_8615_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_d78e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_a882 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_ed3c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_7e32 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_uxn_opcodes_h_l1372_c3_8871 : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_return_output : unsigned(8 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_c5a1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_a19e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_80dc : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_uxn_opcodes_h_l1379_c3_25e0 : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_left : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_8615_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_8615_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_8615_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_8615_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c99_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_692b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4ac1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_279e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1351_l1386_DUPLICATE_a0f7_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_7e32 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_7e32;
     VAR_MUX_uxn_opcodes_h_l1379_c37_8615_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_c5a1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_c5a1;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1379_c37_8615_iffalse := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_a882 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_a882;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_ed3c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_ed3c;
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_d78e := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_d78e;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_80dc := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_80dc;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_left := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_left := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse := t16_high;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_left := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse := t16_low;
     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1371_c11_b1b1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1379_c37_bc63] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_left;
     BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_return_output := BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1368_c11_df5f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1372_c13_5bb4] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output := result.is_ram_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1378_c7_a19e] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_a19e_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_0fa0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l1373_c30_09f9] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_ins;
     sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_x;
     sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_return_output := sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c99 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c99_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4ac1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4ac1_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_279e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_279e_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1355_c6_1f9a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_692b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_692b_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_1f9a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_df5f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_b1b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_0fa0_return_output;
     VAR_MUX_uxn_opcodes_h_l1379_c37_8615_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_bc63_return_output;
     VAR_t16_low_uxn_opcodes_h_l1372_c3_8871 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_5bb4_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_692b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_692b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_279e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_279e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_279e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4ac1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_4ac1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c99_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c99_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c99_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_36cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_a19e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_09f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue := VAR_t16_low_uxn_opcodes_h_l1372_c3_8871;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue := VAR_t16_low_uxn_opcodes_h_l1372_c3_8871;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1371_c7_9acb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_a19e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c7_a19e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;

     -- MUX[uxn_opcodes_h_l1379_c37_8615] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1379_c37_8615_cond <= VAR_MUX_uxn_opcodes_h_l1379_c37_8615_cond;
     MUX_uxn_opcodes_h_l1379_c37_8615_iftrue <= VAR_MUX_uxn_opcodes_h_l1379_c37_8615_iftrue;
     MUX_uxn_opcodes_h_l1379_c37_8615_iffalse <= VAR_MUX_uxn_opcodes_h_l1379_c37_8615_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1379_c37_8615_return_output := MUX_uxn_opcodes_h_l1379_c37_8615_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_a19e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1371_c7_9acb] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_cond;
     t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output := t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_right := VAR_MUX_uxn_opcodes_h_l1379_c37_8615_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1371_c7_9acb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1368_c7_aa69] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1379_c14_6259] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1371_c7_9acb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1368_c7_aa69] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_cond;
     t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output := t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1371_c7_9acb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;

     -- Submodule level 3
     VAR_t16_high_uxn_opcodes_h_l1379_c3_25e0 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_6259_return_output, 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue := VAR_t16_high_uxn_opcodes_h_l1379_c3_25e0;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue := VAR_t16_high_uxn_opcodes_h_l1379_c3_25e0;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1368_c7_aa69] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1368_c7_aa69] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1368_c7_aa69] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_a19e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1378_c7_a19e] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_cond;
     t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output := t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_a19e_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1371_c7_9acb] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_cond;
     t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output := t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1371_c7_9acb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- Submodule level 5
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_9acb_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1368_c7_aa69] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output := result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1368_c7_aa69] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_cond;
     t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output := t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_aa69_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1355_c2_36cc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;

     -- Submodule level 7
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1351_l1386_DUPLICATE_a0f7 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1351_l1386_DUPLICATE_a0f7_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_36cc_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1351_l1386_DUPLICATE_a0f7_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e6e6_uxn_opcodes_h_l1351_l1386_DUPLICATE_a0f7_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
