-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 36
entity nip2_0CLK_1a2ef46d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_1a2ef46d;
architecture arch of nip2_0CLK_1a2ef46d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2174_c6_9304]
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2174_c2_f3fe]
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_ce34]
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2187_c7_f3ff]
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_f3ff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_f3ff]
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_f3ff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_f3ff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_f3ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2187_c7_f3ff]
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_65d3]
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2190_c7_c836]
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_c836]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_c836]
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_c836]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_c836]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_c836]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2190_c7_c836]
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2192_c30_9c1c]
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_09d5]
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2197_c7_0c30]
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_0c30]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_0c30]
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_0c30]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_0c30]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_b856( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_left,
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_right,
BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe
t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe
t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond,
t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue,
t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse,
t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_left,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_right,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff
t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond,
t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue,
t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse,
t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff
t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond,
t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue,
t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse,
t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_left,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_right,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2190_c7_c836
t16_low_MUX_uxn_opcodes_h_l2190_c7_c836 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_cond,
t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue,
t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse,
t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_cond,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2190_c7_c836
t16_high_MUX_uxn_opcodes_h_l2190_c7_c836 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_cond,
t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue,
t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse,
t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c
sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_ins,
sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_x,
sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_y,
sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_left,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_right,
BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30
t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_cond,
t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue,
t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse,
t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_cond,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output,
 t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output,
 t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output,
 t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output,
 t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_return_output,
 t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_return_output,
 sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output,
 t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_14ad : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_db04 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_7e71 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_0ae2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_23cf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_0c30_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_2773 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_303d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_0015_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_2013_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_87ed_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2205_l2170_DUPLICATE_daa5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_14ad := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2184_c3_14ad;
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_7e71 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2188_c3_7e71;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_23cf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2200_c3_23cf;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_db04 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2179_c3_db04;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_2773 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2199_c3_2773;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_0ae2 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2194_c3_0ae2;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse := t16_high;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse := t16_low;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2197_c7_0c30] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_0c30_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_ce34] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_left;
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output := BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_303d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_303d_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_0015 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_0015_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2197_c11_09d5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_2013 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_2013_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2174_c6_9304] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_left;
     BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output := BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_65d3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l2192_c30_9c1c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_ins;
     sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_x;
     sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_return_output := sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_87ed LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_87ed_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2174_c6_9304_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_ce34_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_65d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c11_09d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_2013_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2197_l2187_DUPLICATE_2013_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_87ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_87ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2197_l2187_l2190_DUPLICATE_87ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_0015_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_0015_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_303d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_303d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2174_l2197_l2187_DUPLICATE_303d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2174_c2_f3fe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2197_c7_0c30_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2192_c30_9c1c_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2190_c7_c836] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_cond;
     t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_return_output := t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c7_0c30] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_c836] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2197_c7_0c30] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_cond;
     t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output := t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2197_c7_0c30] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output := result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c7_0c30] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c7_0c30] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2197_c7_0c30_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2187_c7_f3ff] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond;
     t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output := t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_c836] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_return_output := result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_c836] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_f3ff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_c836] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_c836] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2190_c7_c836] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_cond;
     t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_return_output := t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2190_c7_c836_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2187_c7_f3ff] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond;
     t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output := t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_f3ff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_f3ff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output := result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_f3ff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_f3ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2187_c7_f3ff_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2174_c2_f3fe] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;

     -- Submodule level 5
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2205_l2170_DUPLICATE_daa5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2205_l2170_DUPLICATE_daa5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_b856(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2174_c2_f3fe_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2205_l2170_DUPLICATE_daa5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_b856_uxn_opcodes_h_l2205_l2170_DUPLICATE_daa5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
