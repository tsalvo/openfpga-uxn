-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity mul_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_64d180f1;
architecture arch of mul_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1987_c6_49a3]
signal BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1987_c2_3c2f]
signal n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2000_c11_6fe5]
signal BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2000_c7_3139]
signal t8_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2000_c7_3139]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2000_c7_3139]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2000_c7_3139]
signal result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2000_c7_3139]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2000_c7_3139]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2000_c7_3139]
signal n8_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2003_c11_0393]
signal BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2003_c7_52a7]
signal t8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2003_c7_52a7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2003_c7_52a7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2003_c7_52a7]
signal result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2003_c7_52a7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2003_c7_52a7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2003_c7_52a7]
signal n8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2006_c11_7e9f]
signal BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2006_c7_01b1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2006_c7_01b1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2006_c7_01b1]
signal result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2006_c7_01b1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2006_c7_01b1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2006_c7_01b1]
signal n8_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2008_c30_66f0]
signal sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2011_c21_0c42]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_return_output : unsigned(15 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c580( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3
BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_left,
BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_right,
BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output);

-- t8_MUX_uxn_opcodes_h_l1987_c2_3c2f
t8_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f
result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- n8_MUX_uxn_opcodes_h_l1987_c2_3c2f
n8_MUX_uxn_opcodes_h_l1987_c2_3c2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond,
n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue,
n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse,
n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5
BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_left,
BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_right,
BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output);

-- t8_MUX_uxn_opcodes_h_l2000_c7_3139
t8_MUX_uxn_opcodes_h_l2000_c7_3139 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2000_c7_3139_cond,
t8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue,
t8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse,
t8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139
result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139
result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_cond,
result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139
result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139
result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_return_output);

-- n8_MUX_uxn_opcodes_h_l2000_c7_3139
n8_MUX_uxn_opcodes_h_l2000_c7_3139 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2000_c7_3139_cond,
n8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue,
n8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse,
n8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393
BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_left,
BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_right,
BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output);

-- t8_MUX_uxn_opcodes_h_l2003_c7_52a7
t8_MUX_uxn_opcodes_h_l2003_c7_52a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond,
t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue,
t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse,
t8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7
result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7
result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7
result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output);

-- n8_MUX_uxn_opcodes_h_l2003_c7_52a7
n8_MUX_uxn_opcodes_h_l2003_c7_52a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond,
n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue,
n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse,
n8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f
BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_left,
BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_right,
BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1
result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1
result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1
result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output);

-- n8_MUX_uxn_opcodes_h_l2006_c7_01b1
n8_MUX_uxn_opcodes_h_l2006_c7_01b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2006_c7_01b1_cond,
n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue,
n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse,
n8_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0
sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_ins,
sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_x,
sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_y,
sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42 : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output,
 t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output,
 t8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_return_output,
 n8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output,
 t8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output,
 n8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output,
 n8_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output,
 sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1997_c3_a741 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1992_c3_972b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2001_c3_16bb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2010_c3_91e5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l2011_c3_709b : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2003_l1987_l2006_l2000_DUPLICATE_26ae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_372a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_4a0c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_ec82_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2003_l2006_DUPLICATE_aa02_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2015_l1983_DUPLICATE_b688_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1992_c3_972b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1992_c3_972b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2010_c3_91e5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2010_c3_91e5;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1997_c3_a741 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1997_c3_a741;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2001_c3_16bb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2001_c3_16bb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1987_c6_49a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_left;
     BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output := BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2003_l1987_l2006_l2000_DUPLICATE_26ae LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2003_l1987_l2006_l2000_DUPLICATE_26ae_return_output := result.u8_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2006_c11_7e9f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l2008_c30_66f0] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_ins;
     sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_x;
     sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_return_output := sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_ec82 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_ec82_return_output := result.sp_relative_shift;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2011_c21_0c42] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_372a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_372a_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_4a0c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_4a0c_return_output := result.is_stack_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output := result.is_pc_updated;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2003_c11_0393] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_left;
     BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output := BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2000_c11_6fe5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2003_l2006_DUPLICATE_aa02 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2003_l2006_DUPLICATE_aa02_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1987_c6_49a3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2000_c11_6fe5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2003_c11_0393_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2006_c11_7e9f_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l2011_c3_709b := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2011_c21_0c42_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_ec82_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_ec82_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_ec82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_372a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_372a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_372a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_4a0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_4a0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2003_l2006_l2000_DUPLICATE_4a0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2003_l2006_DUPLICATE_aa02_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2003_l2006_DUPLICATE_aa02_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2003_l1987_l2006_l2000_DUPLICATE_26ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2003_l1987_l2006_l2000_DUPLICATE_26ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2003_l1987_l2006_l2000_DUPLICATE_26ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2003_l1987_l2006_l2000_DUPLICATE_26ae_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1987_c2_3c2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2008_c30_66f0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue := VAR_result_u8_value_uxn_opcodes_h_l2011_c3_709b;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2006_c7_01b1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;

     -- n8_MUX[uxn_opcodes_h_l2006_c7_01b1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2006_c7_01b1_cond <= VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_cond;
     n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue;
     n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output := n8_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2003_c7_52a7] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond <= VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond;
     t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue;
     t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output := t8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2006_c7_01b1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2006_c7_01b1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2006_c7_01b1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2006_c7_01b1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2006_c7_01b1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2003_c7_52a7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2003_c7_52a7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2003_c7_52a7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;

     -- n8_MUX[uxn_opcodes_h_l2003_c7_52a7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond <= VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_cond;
     n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue;
     n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output := n8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2003_c7_52a7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;

     -- t8_MUX[uxn_opcodes_h_l2000_c7_3139] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2000_c7_3139_cond <= VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_cond;
     t8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue;
     t8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output := t8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2003_c7_52a7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2003_c7_52a7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;
     -- n8_MUX[uxn_opcodes_h_l2000_c7_3139] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2000_c7_3139_cond <= VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_cond;
     n8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue;
     n8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output := n8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2000_c7_3139] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_return_output := result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;

     -- t8_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2000_c7_3139] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2000_c7_3139] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2000_c7_3139] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2000_c7_3139] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2000_c7_3139_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- n8_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1987_c2_3c2f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2015_l1983_DUPLICATE_b688 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2015_l1983_DUPLICATE_b688_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c580(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1987_c2_3c2f_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2015_l1983_DUPLICATE_b688_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2015_l1983_DUPLICATE_b688_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
