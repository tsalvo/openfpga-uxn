-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity dup_0CLK_a148083c is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_a148083c;
architecture arch of dup_0CLK_a148083c is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2566_c6_bd40]
signal BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2566_c1_04f9]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2566_c2_c565]
signal t8_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2566_c2_c565]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2566_c2_c565]
signal result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2566_c2_c565]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2566_c2_c565]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2566_c2_c565]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2566_c2_c565]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2566_c2_c565]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l2567_c3_75d6[uxn_opcodes_h_l2567_c3_75d6]
signal printf_uxn_opcodes_h_l2567_c3_75d6_uxn_opcodes_h_l2567_c3_75d6_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2572_c11_505c]
signal BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2572_c7_c5a6]
signal t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2572_c7_c5a6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2572_c7_c5a6]
signal result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2572_c7_c5a6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2572_c7_c5a6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2572_c7_c5a6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2572_c7_c5a6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2572_c7_c5a6]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2575_c11_29fc]
signal BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2575_c7_3bf4]
signal t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2575_c7_3bf4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2575_c7_3bf4]
signal result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2575_c7_3bf4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2575_c7_3bf4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2575_c7_3bf4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2575_c7_3bf4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(7 downto 0);

-- result_is_stack_read_MUX[uxn_opcodes_h_l2575_c7_3bf4]
signal result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(0 downto 0);
signal result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2579_c32_3d45]
signal BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2579_c32_7579]
signal BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2579_c32_49bd]
signal MUX_uxn_opcodes_h_l2579_c32_49bd_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2579_c32_49bd_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2579_c32_49bd_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2579_c32_49bd_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2581_c11_0ee2]
signal BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2581_c7_aac6]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2581_c7_aac6]
signal result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2581_c7_aac6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2581_c7_aac6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2581_c7_aac6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2587_c11_b1ed]
signal BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2587_c7_7d62]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2587_c7_7d62]
signal result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2587_c7_7d62]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2587_c7_7d62]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2591_c11_06d2]
signal BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2591_c7_2394]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2591_c7_2394]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e56b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_sp_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_stack_read := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40
BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_left,
BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_right,
BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_return_output);

-- t8_MUX_uxn_opcodes_h_l2566_c2_c565
t8_MUX_uxn_opcodes_h_l2566_c2_c565 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2566_c2_c565_cond,
t8_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue,
t8_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse,
t8_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565
result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565
result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_cond,
result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565
result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565
result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565
result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565
result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

-- printf_uxn_opcodes_h_l2567_c3_75d6_uxn_opcodes_h_l2567_c3_75d6
printf_uxn_opcodes_h_l2567_c3_75d6_uxn_opcodes_h_l2567_c3_75d6 : entity work.printf_uxn_opcodes_h_l2567_c3_75d6_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2567_c3_75d6_uxn_opcodes_h_l2567_c3_75d6_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c
BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_left,
BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_right,
BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output);

-- t8_MUX_uxn_opcodes_h_l2572_c7_c5a6
t8_MUX_uxn_opcodes_h_l2572_c7_c5a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond,
t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue,
t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse,
t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6
result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6
result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond,
result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6
result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6
result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6
result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc
BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_left,
BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_right,
BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output);

-- t8_MUX_uxn_opcodes_h_l2575_c7_3bf4
t8_MUX_uxn_opcodes_h_l2575_c7_3bf4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond,
t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue,
t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse,
t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4
result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4
result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond,
result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4
result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4
result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4
result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output);

-- result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4
result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond,
result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue,
result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse,
result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45
BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_left,
BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_right,
BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579
BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_left,
BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_right,
BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_return_output);

-- MUX_uxn_opcodes_h_l2579_c32_49bd
MUX_uxn_opcodes_h_l2579_c32_49bd : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2579_c32_49bd_cond,
MUX_uxn_opcodes_h_l2579_c32_49bd_iftrue,
MUX_uxn_opcodes_h_l2579_c32_49bd_iffalse,
MUX_uxn_opcodes_h_l2579_c32_49bd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2
BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_left,
BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_right,
BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6
result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6
result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_cond,
result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6
result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6
result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed
BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_left,
BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_right,
BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62
result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_cond,
result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62
result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62
result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2
BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_left,
BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_right,
BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394
result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394
result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_return_output,
 t8_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output,
 t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output,
 t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output,
 result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_return_output,
 MUX_uxn_opcodes_h_l2579_c32_49bd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2569_c3_a80a : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2567_c3_75d6_uxn_opcodes_h_l2567_c3_75d6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2573_c3_18e1 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2584_c3_df13 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2588_c3_0224 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2566_l2581_l2572_DUPLICATE_0ae5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2587_l2575_l2566_l2572_DUPLICATE_4557_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2575_l2566_l2572_DUPLICATE_7d9d_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2566_l2591_l2587_l2575_l2572_DUPLICATE_8f03_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2591_l2587_l2581_l2575_l2572_DUPLICATE_0ec3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2575_l2572_DUPLICATE_d9b8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2587_l2575_DUPLICATE_787e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l2596_l2562_DUPLICATE_70a5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2573_c3_18e1 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2573_c3_18e1;
     VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_iftrue := signed(std_logic_vector(resize(to_unsigned(2, 2), 8)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_right := to_unsigned(2, 2);
     VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2569_c3_a80a := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2569_c3_a80a;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_iffalse := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2584_c3_df13 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2584_c3_df13;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_right := to_unsigned(128, 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2588_c3_0224 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2588_c3_0224;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue := VAR_previous_stack_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue := t8;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2575_c11_29fc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_left;
     BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output := BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2575_l2572_DUPLICATE_d9b8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2575_l2572_DUPLICATE_d9b8_return_output := result.is_stack_read;

     -- BIN_OP_EQ[uxn_opcodes_h_l2581_c11_0ee2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2566_c6_bd40] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_left;
     BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output := BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2566_l2581_l2572_DUPLICATE_0ae5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2566_l2581_l2572_DUPLICATE_0ae5_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2591_c11_06d2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2587_l2575_DUPLICATE_787e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2587_l2575_DUPLICATE_787e_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2566_l2591_l2587_l2575_l2572_DUPLICATE_8f03 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2566_l2591_l2587_l2575_l2572_DUPLICATE_8f03_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2572_c11_505c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2587_c11_b1ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2587_l2575_l2566_l2572_DUPLICATE_4557 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2587_l2575_l2566_l2572_DUPLICATE_4557_return_output := result.stack_value;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2575_l2566_l2572_DUPLICATE_7d9d LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2575_l2566_l2572_DUPLICATE_7d9d_return_output := result.sp_relative_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l2579_c32_3d45] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_left;
     BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_return_output := BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2591_l2587_l2581_l2575_l2572_DUPLICATE_0ec3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2591_l2587_l2581_l2575_l2572_DUPLICATE_0ec3_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2579_c32_3d45_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2566_c6_bd40_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2572_c11_505c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2575_c11_29fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2581_c11_0ee2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2587_c11_b1ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2591_c11_06d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2575_l2566_l2572_DUPLICATE_7d9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2575_l2566_l2572_DUPLICATE_7d9d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2575_l2566_l2572_DUPLICATE_7d9d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2591_l2587_l2581_l2575_l2572_DUPLICATE_0ec3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2591_l2587_l2581_l2575_l2572_DUPLICATE_0ec3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2591_l2587_l2581_l2575_l2572_DUPLICATE_0ec3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2591_l2587_l2581_l2575_l2572_DUPLICATE_0ec3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2591_l2587_l2581_l2575_l2572_DUPLICATE_0ec3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2566_l2581_l2572_DUPLICATE_0ae5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2566_l2581_l2572_DUPLICATE_0ae5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2566_l2581_l2572_DUPLICATE_0ae5_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2575_l2572_DUPLICATE_d9b8_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_read_d41d_uxn_opcodes_h_l2575_l2572_DUPLICATE_d9b8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2566_l2591_l2587_l2575_l2572_DUPLICATE_8f03_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2566_l2591_l2587_l2575_l2572_DUPLICATE_8f03_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2566_l2591_l2587_l2575_l2572_DUPLICATE_8f03_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2566_l2591_l2587_l2575_l2572_DUPLICATE_8f03_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2566_l2591_l2587_l2575_l2572_DUPLICATE_8f03_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2587_l2575_DUPLICATE_787e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2587_l2575_DUPLICATE_787e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2587_l2575_l2566_l2572_DUPLICATE_4557_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2587_l2575_l2566_l2572_DUPLICATE_4557_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2587_l2575_l2566_l2572_DUPLICATE_4557_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2587_l2575_l2566_l2572_DUPLICATE_4557_return_output;
     -- BIN_OP_GT[uxn_opcodes_h_l2579_c32_7579] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_left;
     BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_return_output := BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2575_c7_3bf4] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2566_c1_04f9] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2591_c7_2394] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2581_c7_aac6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2575_c7_3bf4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond <= VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond;
     t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue;
     t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output := t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2587_c7_7d62] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output := result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2587_c7_7d62] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2591_c7_2394] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2579_c32_7579_return_output;
     VAR_printf_uxn_opcodes_h_l2567_c3_75d6_uxn_opcodes_h_l2567_c3_75d6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2566_c1_04f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2591_c7_2394_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2591_c7_2394_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;
     -- t8_MUX[uxn_opcodes_h_l2572_c7_c5a6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond;
     t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue;
     t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output := t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2575_c7_3bf4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;

     -- MUX[uxn_opcodes_h_l2579_c32_49bd] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2579_c32_49bd_cond <= VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_cond;
     MUX_uxn_opcodes_h_l2579_c32_49bd_iftrue <= VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_iftrue;
     MUX_uxn_opcodes_h_l2579_c32_49bd_iffalse <= VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_return_output := MUX_uxn_opcodes_h_l2579_c32_49bd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2587_c7_7d62] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2581_c7_aac6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2581_c7_aac6] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output := result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2587_c7_7d62] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output;

     -- printf_uxn_opcodes_h_l2567_c3_75d6[uxn_opcodes_h_l2567_c3_75d6] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2567_c3_75d6_uxn_opcodes_h_l2567_c3_75d6_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2567_c3_75d6_uxn_opcodes_h_l2567_c3_75d6_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2572_c7_c5a6] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue := VAR_MUX_uxn_opcodes_h_l2579_c32_49bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse := VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2587_c7_7d62_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2575_c7_3bf4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2575_c7_3bf4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2581_c7_aac6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2575_c7_3bf4] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output := result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;

     -- t8_MUX[uxn_opcodes_h_l2566_c2_c565] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2566_c2_c565_cond <= VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_cond;
     t8_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue;
     t8_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_return_output := t8_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;

     -- result_is_stack_read_MUX[uxn_opcodes_h_l2566_c2_c565] LATENCY=0
     -- Inputs
     result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_cond <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_cond;
     result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue;
     result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse <= VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse;
     -- Outputs
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_return_output := result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2572_c7_c5a6] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2581_c7_aac6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2581_c7_aac6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2575_c7_3bf4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2572_c7_c5a6] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output := result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2572_c7_c5a6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2575_c7_3bf4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2572_c7_c5a6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2566_c2_c565] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2575_c7_3bf4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2566_c2_c565] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2572_c7_c5a6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2566_c2_c565] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_return_output := result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2572_c7_c5a6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2566_c2_c565] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2572_c7_c5a6_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2566_c2_c565] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2566_c2_c565] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l2596_l2562_DUPLICATE_70a5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l2596_l2562_DUPLICATE_70a5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e56b(
     result,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2566_c2_c565_return_output,
     VAR_result_is_stack_read_MUX_uxn_opcodes_h_l2566_c2_c565_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l2596_l2562_DUPLICATE_70a5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e56b_uxn_opcodes_h_l2596_l2562_DUPLICATE_70a5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
