-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity nip2_0CLK_b2fbb329 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_b2fbb329;
architecture arch of nip2_0CLK_b2fbb329 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2137_c6_950f]
signal BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2137_c2_fe47]
signal t16_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2137_c2_fe47]
signal result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2137_c2_fe47]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2137_c2_fe47]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2137_c2_fe47]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2137_c2_fe47]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2144_c11_e190]
signal BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2144_c7_3e53]
signal t16_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2144_c7_3e53]
signal result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2144_c7_3e53]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2144_c7_3e53]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2144_c7_3e53]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2144_c7_3e53]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2147_c11_b661]
signal BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2147_c7_3e68]
signal t16_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2147_c7_3e68]
signal result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2147_c7_3e68]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2147_c7_3e68]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2147_c7_3e68]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2147_c7_3e68]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : signed(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2149_c3_7cf4]
signal CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2151_c11_f3cb]
signal BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2151_c7_661e]
signal t16_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2151_c7_661e]
signal result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2151_c7_661e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2151_c7_661e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2151_c7_661e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2151_c7_661e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : signed(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2152_c3_af1d]
signal BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2154_c30_39ce]
signal sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2159_c11_fb5a]
signal BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2159_c7_8df0]
signal result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2159_c7_8df0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2159_c7_8df0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2159_c7_8df0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2159_c7_8df0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : signed(3 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l2162_c31_6a85]
signal CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2164_c11_bb7f]
signal BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2164_c7_3d46]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2164_c7_3d46]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f
BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_left,
BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_right,
BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output);

-- t16_MUX_uxn_opcodes_h_l2137_c2_fe47
t16_MUX_uxn_opcodes_h_l2137_c2_fe47 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2137_c2_fe47_cond,
t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue,
t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse,
t16_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47
result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_cond,
result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47
result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47
result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47
result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190
BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_left,
BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_right,
BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output);

-- t16_MUX_uxn_opcodes_h_l2144_c7_3e53
t16_MUX_uxn_opcodes_h_l2144_c7_3e53 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2144_c7_3e53_cond,
t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue,
t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse,
t16_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53
result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_cond,
result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661
BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_left,
BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_right,
BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output);

-- t16_MUX_uxn_opcodes_h_l2147_c7_3e68
t16_MUX_uxn_opcodes_h_l2147_c7_3e68 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2147_c7_3e68_cond,
t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue,
t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse,
t16_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68
result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_cond,
result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4
CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_x,
CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb
BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_left,
BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_right,
BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output);

-- t16_MUX_uxn_opcodes_h_l2151_c7_661e
t16_MUX_uxn_opcodes_h_l2151_c7_661e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2151_c7_661e_cond,
t16_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue,
t16_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse,
t16_MUX_uxn_opcodes_h_l2151_c7_661e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e
result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d
BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_left,
BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_right,
BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce
sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_ins,
sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_x,
sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_y,
sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a
BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_left,
BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_right,
BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0
result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output);

-- CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85
CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_x,
CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f
BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_left,
BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_right,
BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46
result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46
result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output,
 t16_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output,
 t16_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output,
 t16_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output,
 CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output,
 t16_MUX_uxn_opcodes_h_l2151_c7_661e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_return_output,
 sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output,
 CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2141_c3_80b9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2145_c3_d1f4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2156_c3_ff4c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2157_c21_98c3_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2161_c3_d9a5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2160_c3_d93b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2162_c21_4f81_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_4bf8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2144_l2137_l2164_l2147_l2159_DUPLICATE_c12d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_efb4_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2151_l2144_l2164_l2147_l2159_DUPLICATE_ffef_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2148_l2152_DUPLICATE_c6d9_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2147_l2159_DUPLICATE_ae4b_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2169_l2133_DUPLICATE_c60b_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2161_c3_d9a5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2161_c3_d9a5;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2156_c3_ff4c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2156_c3_ff4c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2141_c3_80b9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2141_c3_80b9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2145_c3_d1f4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2145_c3_d1f4;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_y := resize(to_signed(-2, 3), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2160_c3_d93b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2160_c3_d93b;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_left := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_x := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse := t16;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_4bf8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_4bf8_return_output := result.u8_value;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2148_l2152_DUPLICATE_c6d9 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2148_l2152_DUPLICATE_c6d9_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2151_c11_f3cb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2144_c11_e190] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_left;
     BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output := BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l2162_c31_6a85] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_x <= VAR_CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_return_output := CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2144_l2137_l2164_l2147_l2159_DUPLICATE_c12d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2144_l2137_l2164_l2147_l2159_DUPLICATE_c12d_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2159_c11_fb5a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2164_c11_bb7f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2147_l2159_DUPLICATE_ae4b LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2147_l2159_DUPLICATE_ae4b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2137_c6_950f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2147_c11_b661] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_left;
     BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output := BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2151_l2144_l2164_l2147_l2159_DUPLICATE_ffef LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2151_l2144_l2164_l2147_l2159_DUPLICATE_ffef_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l2154_c30_39ce] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_ins;
     sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_x;
     sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_return_output := sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_efb4 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_efb4_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2137_c6_950f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_e190_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_b661_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_f3cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_fb5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2164_c11_bb7f_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2148_l2152_DUPLICATE_c6d9_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2148_l2152_DUPLICATE_c6d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_efb4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_efb4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_efb4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_efb4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2151_l2144_l2164_l2147_l2159_DUPLICATE_ffef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2151_l2144_l2164_l2147_l2159_DUPLICATE_ffef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2151_l2144_l2164_l2147_l2159_DUPLICATE_ffef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2151_l2144_l2164_l2147_l2159_DUPLICATE_ffef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2151_l2144_l2164_l2147_l2159_DUPLICATE_ffef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2144_l2137_l2164_l2147_l2159_DUPLICATE_c12d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2144_l2137_l2164_l2147_l2159_DUPLICATE_c12d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2144_l2137_l2164_l2147_l2159_DUPLICATE_c12d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2144_l2137_l2164_l2147_l2159_DUPLICATE_c12d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2144_l2137_l2164_l2147_l2159_DUPLICATE_c12d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2147_l2159_DUPLICATE_ae4b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2147_l2159_DUPLICATE_ae4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_4bf8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_4bf8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_4bf8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2147_l2137_l2159_l2144_DUPLICATE_4bf8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2154_c30_39ce_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2164_c7_3d46] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2159_c7_8df0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2152_c3_af1d] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_left;
     BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_return_output := BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2164_c7_3d46] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2162_c21_4f81] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2162_c21_4f81_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l2162_c31_6a85_return_output);

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2159_c7_8df0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2149_c3_7cf4] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_return_output := CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2162_c21_4f81_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2149_c3_7cf4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2164_c7_3d46_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2151_c7_661e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2159_c7_8df0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2159_c7_8df0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2157_c21_98c3] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2157_c21_98c3_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l2152_c3_af1d_return_output);

     -- t16_MUX[uxn_opcodes_h_l2151_c7_661e] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2151_c7_661e_cond <= VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_cond;
     t16_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue;
     t16_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_return_output := t16_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2159_c7_8df0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2151_c7_661e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2157_c21_98c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2159_c7_8df0_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2151_c7_661e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2151_c7_661e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2147_c7_3e68] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2147_c7_3e68] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;

     -- t16_MUX[uxn_opcodes_h_l2147_c7_3e68] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2147_c7_3e68_cond <= VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_cond;
     t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue;
     t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output := t16_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2151_c7_661e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2151_c7_661e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;
     -- t16_MUX[uxn_opcodes_h_l2144_c7_3e53] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2144_c7_3e53_cond <= VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_cond;
     t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue;
     t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output := t16_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2144_c7_3e53] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2144_c7_3e53] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2147_c7_3e68] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2147_c7_3e68] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2147_c7_3e68] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output := result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2147_c7_3e68_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2137_c2_fe47] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output;

     -- t16_MUX[uxn_opcodes_h_l2137_c2_fe47] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2137_c2_fe47_cond <= VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_cond;
     t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue;
     t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output := t16_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2137_c2_fe47] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2144_c7_3e53] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2144_c7_3e53] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2144_c7_3e53] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output := result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2144_c7_3e53_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2137_c2_fe47] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2137_c2_fe47] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2137_c2_fe47] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output := result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2169_l2133_DUPLICATE_c60b LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2169_l2133_DUPLICATE_c60b_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2137_c2_fe47_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2169_l2133_DUPLICATE_c60b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2169_l2133_DUPLICATE_c60b_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
