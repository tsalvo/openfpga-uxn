-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_0490]
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal l8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal t8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2639_c2_76b6]
signal n8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_5001]
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2652_c7_8c06]
signal l8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2652_c7_8c06]
signal t8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_8c06]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_8c06]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_8c06]
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_8c06]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_8c06]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2652_c7_8c06]
signal n8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_4edf]
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2655_c7_93d6]
signal l8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2655_c7_93d6]
signal t8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_93d6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_93d6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_93d6]
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_93d6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_93d6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2655_c7_93d6]
signal n8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_6693]
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2659_c7_9d5a]
signal l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_9d5a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_9d5a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_9d5a]
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_9d5a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_9d5a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2659_c7_9d5a]
signal n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2661_c30_708d]
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_4dcb]
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2666_c7_5ffd]
signal l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_5ffd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_5ffd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_5ffd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_5ffd]
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_6b34]
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_6cbf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_6cbf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_6cbf]
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_71f0( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_index_flipped := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_left,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_right,
BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output);

-- l8_MUX_uxn_opcodes_h_l2639_c2_76b6
l8_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
l8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- t8_MUX_uxn_opcodes_h_l2639_c2_76b6
t8_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
t8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- n8_MUX_uxn_opcodes_h_l2639_c2_76b6
n8_MUX_uxn_opcodes_h_l2639_c2_76b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond,
n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue,
n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse,
n8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_left,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_right,
BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output);

-- l8_MUX_uxn_opcodes_h_l2652_c7_8c06
l8_MUX_uxn_opcodes_h_l2652_c7_8c06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond,
l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue,
l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse,
l8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output);

-- t8_MUX_uxn_opcodes_h_l2652_c7_8c06
t8_MUX_uxn_opcodes_h_l2652_c7_8c06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond,
t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue,
t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse,
t8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_cond,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output);

-- n8_MUX_uxn_opcodes_h_l2652_c7_8c06
n8_MUX_uxn_opcodes_h_l2652_c7_8c06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond,
n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue,
n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse,
n8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_left,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_right,
BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output);

-- l8_MUX_uxn_opcodes_h_l2655_c7_93d6
l8_MUX_uxn_opcodes_h_l2655_c7_93d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond,
l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue,
l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse,
l8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output);

-- t8_MUX_uxn_opcodes_h_l2655_c7_93d6
t8_MUX_uxn_opcodes_h_l2655_c7_93d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond,
t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue,
t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse,
t8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output);

-- n8_MUX_uxn_opcodes_h_l2655_c7_93d6
n8_MUX_uxn_opcodes_h_l2655_c7_93d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond,
n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue,
n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse,
n8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_left,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_right,
BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output);

-- l8_MUX_uxn_opcodes_h_l2659_c7_9d5a
l8_MUX_uxn_opcodes_h_l2659_c7_9d5a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond,
l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue,
l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse,
l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output);

-- n8_MUX_uxn_opcodes_h_l2659_c7_9d5a
n8_MUX_uxn_opcodes_h_l2659_c7_9d5a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond,
n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue,
n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse,
n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2661_c30_708d
sp_relative_shift_uxn_opcodes_h_l2661_c30_708d : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_ins,
sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_x,
sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_y,
sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_left,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_right,
BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output);

-- l8_MUX_uxn_opcodes_h_l2666_c7_5ffd
l8_MUX_uxn_opcodes_h_l2666_c7_5ffd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond,
l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue,
l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse,
l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_left,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_right,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output,
 l8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 t8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 n8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output,
 l8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output,
 t8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output,
 n8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output,
 l8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output,
 t8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output,
 n8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output,
 l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output,
 n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output,
 sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output,
 l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_6b76 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_716f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_e16b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_bf32 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_2f19 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_797b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_d96f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_3046 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_6cbf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2672_l2639_l2652_DUPLICATE_e73c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_429c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2652_l2666_DUPLICATE_18cb_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_69ef_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2678_l2635_DUPLICATE_955a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_6b76 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2644_c3_6b76;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_3046 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_3046;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_2f19 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2663_c3_2f19;
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_e16b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2653_c3_e16b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_bf32 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2656_c3_bf32;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_716f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2649_c3_716f;
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_d96f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2668_c3_d96f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_797b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2669_c3_797b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_right := to_unsigned(5, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse := t8;
     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_429c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_429c_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2659_c11_6693] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_left;
     BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output := BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2652_c11_5001] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_left;
     BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output := BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2672_c7_6cbf] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_6cbf_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2672_l2639_l2652_DUPLICATE_e73c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2672_l2639_l2652_DUPLICATE_e73c_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_6b34] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_left;
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output := BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2652_l2666_DUPLICATE_18cb LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2652_l2666_DUPLICATE_18cb_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2666_c11_4dcb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2661_c30_708d] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_ins;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_x;
     sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_return_output := sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2655_c11_4edf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_left;
     BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output := BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_69ef LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_69ef_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2639_c6_0490] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_left;
     BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output := BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c6_0490_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2652_c11_5001_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2655_c11_4edf_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2659_c11_6693_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2666_c11_4dcb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_6b34_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2652_l2666_DUPLICATE_18cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2652_l2666_DUPLICATE_18cb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2655_l2652_l2666_DUPLICATE_18cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_69ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_69ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_69ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_69ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2672_l2666_l2659_l2655_l2652_DUPLICATE_69ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_429c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_429c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2655_l2659_l2652_DUPLICATE_429c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2672_l2639_l2652_DUPLICATE_e73c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2672_l2639_l2652_DUPLICATE_e73c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2672_l2639_l2652_DUPLICATE_e73c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2655_l2672_l2639_l2652_DUPLICATE_e73c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2639_c2_76b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2672_c7_6cbf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2661_c30_708d_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2666_c7_5ffd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;

     -- t8_MUX[uxn_opcodes_h_l2655_c7_93d6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond;
     t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue;
     t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output := t8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_6cbf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output := result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- l8_MUX[uxn_opcodes_h_l2666_c7_5ffd] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond;
     l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue;
     l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output := l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_6cbf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output;

     -- n8_MUX[uxn_opcodes_h_l2659_c7_9d5a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond;
     n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue;
     n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output := n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2659_c7_9d5a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_6cbf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_6cbf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2655_c7_93d6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;

     -- t8_MUX[uxn_opcodes_h_l2652_c7_8c06] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond;
     t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue;
     t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output := t8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2666_c7_5ffd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2659_c7_9d5a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2666_c7_5ffd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output := result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2666_c7_5ffd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;

     -- n8_MUX[uxn_opcodes_h_l2655_c7_93d6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond;
     n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue;
     n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output := n8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;

     -- l8_MUX[uxn_opcodes_h_l2659_c7_9d5a] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond;
     l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue;
     l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output := l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2666_c7_5ffd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2652_c7_8c06] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;

     -- l8_MUX[uxn_opcodes_h_l2655_c7_93d6] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_cond;
     l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue;
     l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output := l8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2655_c7_93d6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2659_c7_9d5a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := t8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2652_c7_8c06] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond;
     n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue;
     n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output := n8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2659_c7_9d5a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2659_c7_9d5a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2659_c7_9d5a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2655_c7_93d6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2652_c7_8c06] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2655_c7_93d6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;

     -- n8_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := n8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- l8_MUX[uxn_opcodes_h_l2652_c7_8c06] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_cond;
     l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue;
     l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output := l8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2655_c7_93d6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2655_c7_93d6_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2652_c7_8c06] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2652_c7_8c06] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2652_c7_8c06] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output := result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;

     -- l8_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := l8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2652_c7_8c06_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c2_76b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2678_l2635_DUPLICATE_955a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2678_l2635_DUPLICATE_955a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_71f0(
     result,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c2_76b6_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2678_l2635_DUPLICATE_955a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_71f0_uxn_opcodes_h_l2678_l2635_DUPLICATE_955a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
