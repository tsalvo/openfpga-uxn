-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity inc2_0CLK_180c5210 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_180c5210;
architecture arch of inc2_0CLK_180c5210 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1356_c6_36ec]
signal BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1356_c2_1f79]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1369_c11_3c7d]
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1369_c7_28da]
signal t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1369_c7_28da]
signal t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1369_c7_28da]
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1369_c7_28da]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1369_c7_28da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1369_c7_28da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1369_c7_28da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1372_c11_9a77]
signal BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1372_c7_6a67]
signal t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1372_c7_6a67]
signal t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1372_c7_6a67]
signal result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1372_c7_6a67]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1372_c7_6a67]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1372_c7_6a67]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1372_c7_6a67]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1373_c13_ad7b]
signal BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_return_output : unsigned(8 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1374_c30_6072]
signal sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1379_c11_83c7]
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1379_c7_b8d9]
signal t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1379_c7_b8d9]
signal result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1379_c7_b8d9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1379_c7_b8d9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1379_c7_b8d9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1380_c37_c61a]
signal BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1380_c37_6643]
signal MUX_uxn_opcodes_h_l1380_c37_6643_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1380_c37_6643_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1380_c37_6643_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1380_c37_6643_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1380_c14_e9ef]
signal BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_243c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec
BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_left,
BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_right,
BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79
t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79
t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79
result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79
result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79
result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79
result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79
result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79
result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79
result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d
BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_left,
BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_right,
BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1369_c7_28da
t16_low_MUX_uxn_opcodes_h_l1369_c7_28da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_cond,
t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue,
t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse,
t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1369_c7_28da
t16_high_MUX_uxn_opcodes_h_l1369_c7_28da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_cond,
t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue,
t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse,
t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_cond,
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77
BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_left,
BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_right,
BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67
t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_cond,
t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue,
t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse,
t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67
t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_cond,
t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue,
t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse,
t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67
result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_cond,
result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67
result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67
result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67
result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b
BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_left,
BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_right,
BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1374_c30_6072
sp_relative_shift_uxn_opcodes_h_l1374_c30_6072 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_ins,
sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_x,
sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_y,
sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7
BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_left,
BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_right,
BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9
t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond,
t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue,
t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse,
t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9
result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9
result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a
BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_left,
BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_right,
BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_return_output);

-- MUX_uxn_opcodes_h_l1380_c37_6643
MUX_uxn_opcodes_h_l1380_c37_6643 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1380_c37_6643_cond,
MUX_uxn_opcodes_h_l1380_c37_6643_iftrue,
MUX_uxn_opcodes_h_l1380_c37_6643_iffalse,
MUX_uxn_opcodes_h_l1380_c37_6643_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef
BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_left,
BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_right,
BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output,
 t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output,
 t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_return_output,
 t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output,
 t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output,
 t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output,
 t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_return_output,
 MUX_uxn_opcodes_h_l1380_c37_6643_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1366_c3_a346 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1361_c3_2fc2 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1370_c3_f4d2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_uxn_opcodes_h_l1373_c3_6256 : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1376_c3_f6e1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_return_output : unsigned(8 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_uxn_opcodes_h_l1380_c3_1f69 : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1381_c3_8d64 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1382_c3_6e62 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1379_c7_b8d9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_left : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1380_c37_6643_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1380_c37_6643_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1380_c37_6643_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1380_c37_6643_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1356_l1379_l1369_DUPLICATE_023c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1372_l1369_DUPLICATE_7cc6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1379_l1369_DUPLICATE_98e5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1372_l1379_l1369_DUPLICATE_54f3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1352_l1387_DUPLICATE_9b15_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l1380_c37_6643_iffalse := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1382_c3_6e62 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1382_c3_6e62;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1381_c3_8d64 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1381_c3_8d64;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1366_c3_a346 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1366_c3_a346;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1370_c3_f4d2 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1370_c3_f4d2;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_right := to_unsigned(3, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1376_c3_f6e1 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1376_c3_f6e1;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1361_c3_2fc2 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1361_c3_2fc2;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1380_c37_6643_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_left := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_left := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse := t16_high;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_left := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse := t16_low;
     -- sp_relative_shift[uxn_opcodes_h_l1374_c30_6072] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_ins;
     sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_x;
     sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_return_output := sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1369_c11_3c7d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1372_l1369_DUPLICATE_7cc6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1372_l1369_DUPLICATE_7cc6_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1379_l1369_DUPLICATE_98e5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1379_l1369_DUPLICATE_98e5_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1379_c7_b8d9] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1379_c7_b8d9_return_output := result.stack_address_sp_offset;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1373_c13_ad7b] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1380_c37_c61a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1356_l1379_l1369_DUPLICATE_023c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1356_l1379_l1369_DUPLICATE_023c_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1372_l1379_l1369_DUPLICATE_54f3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1372_l1379_l1369_DUPLICATE_54f3_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1379_c11_83c7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_left;
     BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output := BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output := result.is_stack_index_flipped;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1372_c11_9a77] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_left;
     BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output := BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1356_c6_36ec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_left;
     BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output := BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1356_c6_36ec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1369_c11_3c7d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1372_c11_9a77_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c11_83c7_return_output;
     VAR_MUX_uxn_opcodes_h_l1380_c37_6643_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1380_c37_c61a_return_output;
     VAR_t16_low_uxn_opcodes_h_l1373_c3_6256 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1373_c13_ad7b_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1379_l1369_DUPLICATE_98e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1379_l1369_DUPLICATE_98e5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1372_l1379_l1369_DUPLICATE_54f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1372_l1379_l1369_DUPLICATE_54f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1372_l1379_l1369_DUPLICATE_54f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1372_l1369_DUPLICATE_7cc6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1372_l1369_DUPLICATE_7cc6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1356_l1379_l1369_DUPLICATE_023c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1356_l1379_l1369_DUPLICATE_023c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1356_l1379_l1369_DUPLICATE_023c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1356_c2_1f79_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1379_c7_b8d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1374_c30_6072_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue := VAR_t16_low_uxn_opcodes_h_l1373_c3_6256;
     VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue := VAR_t16_low_uxn_opcodes_h_l1373_c3_6256;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1379_c7_b8d9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;

     -- MUX[uxn_opcodes_h_l1380_c37_6643] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1380_c37_6643_cond <= VAR_MUX_uxn_opcodes_h_l1380_c37_6643_cond;
     MUX_uxn_opcodes_h_l1380_c37_6643_iftrue <= VAR_MUX_uxn_opcodes_h_l1380_c37_6643_iftrue;
     MUX_uxn_opcodes_h_l1380_c37_6643_iffalse <= VAR_MUX_uxn_opcodes_h_l1380_c37_6643_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1380_c37_6643_return_output := MUX_uxn_opcodes_h_l1380_c37_6643_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1372_c7_6a67] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_cond;
     t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output := t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1379_c7_b8d9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1379_c7_b8d9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1372_c7_6a67] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_right := VAR_MUX_uxn_opcodes_h_l1380_c37_6643_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1372_c7_6a67] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1369_c7_28da] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_cond;
     t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_return_output := t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1369_c7_28da] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1372_c7_6a67] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1380_c14_e9ef] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1372_c7_6a67] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;

     -- Submodule level 3
     VAR_t16_high_uxn_opcodes_h_l1380_c3_1f69 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1380_c14_e9ef_return_output, 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue := VAR_t16_high_uxn_opcodes_h_l1380_c3_1f69;
     VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue := VAR_t16_high_uxn_opcodes_h_l1380_c3_1f69;
     -- result_u8_value_MUX[uxn_opcodes_h_l1379_c7_b8d9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1369_c7_28da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1369_c7_28da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1379_c7_b8d9] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_cond;
     t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output := t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1369_c7_28da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1379_c7_b8d9_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1372_c7_6a67] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output := result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1372_c7_6a67] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_cond;
     t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output := t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;

     -- Submodule level 5
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1372_c7_6a67_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1369_c7_28da] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_return_output := result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1369_c7_28da] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_cond;
     t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_return_output := t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1369_c7_28da_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1356_c2_1f79] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output := result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;

     -- Submodule level 7
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1352_l1387_DUPLICATE_9b15 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1352_l1387_DUPLICATE_9b15_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_243c(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1356_c2_1f79_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1352_l1387_DUPLICATE_9b15_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_243c_uxn_opcodes_h_l1352_l1387_DUPLICATE_9b15_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
