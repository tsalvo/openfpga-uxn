-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity sta_0CLK_9a874500 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sta_0CLK_9a874500;
architecture arch of sta_0CLK_9a874500 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2258_c6_d2c6]
signal BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2258_c2_8d8f]
signal n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2258_c2_8d8f]
signal t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2258_c2_8d8f]
signal result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2258_c2_8d8f]
signal result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2258_c2_8d8f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2258_c2_8d8f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2258_c2_8d8f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2258_c2_8d8f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2265_c11_d60e]
signal BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2265_c7_2b90]
signal n8_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2265_c7_2b90]
signal t16_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2265_c7_2b90]
signal result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2265_c7_2b90]
signal result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2265_c7_2b90]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2265_c7_2b90]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2265_c7_2b90]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2265_c7_2b90]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2268_c11_cb11]
signal BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2268_c7_fe9f]
signal n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2268_c7_fe9f]
signal t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2268_c7_fe9f]
signal result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2268_c7_fe9f]
signal result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2268_c7_fe9f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2268_c7_fe9f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2268_c7_fe9f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2268_c7_fe9f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(0 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2270_c3_051f]
signal CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2273_c11_2429]
signal BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2273_c7_1ce9]
signal n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2273_c7_1ce9]
signal t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2273_c7_1ce9]
signal result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2273_c7_1ce9]
signal result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2273_c7_1ce9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2273_c7_1ce9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2273_c7_1ce9]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(0 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2274_c3_b7ee]
signal BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2276_c11_43e1]
signal BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2276_c7_531c]
signal n8_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2276_c7_531c]
signal result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2276_c7_531c]
signal result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2276_c7_531c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2276_c7_531c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2276_c7_531c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2279_c30_c336]
signal sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2284_c11_d771]
signal BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2284_c7_ea4f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2284_c7_ea4f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2284_c7_ea4f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_7ccb( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_ram_write := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6
BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_left,
BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_right,
BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output);

-- n8_MUX_uxn_opcodes_h_l2258_c2_8d8f
n8_MUX_uxn_opcodes_h_l2258_c2_8d8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond,
n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue,
n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse,
n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

-- t16_MUX_uxn_opcodes_h_l2258_c2_8d8f
t16_MUX_uxn_opcodes_h_l2258_c2_8d8f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond,
t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue,
t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse,
t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f
result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond,
result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f
result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f
result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f
result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e
BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_left,
BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_right,
BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output);

-- n8_MUX_uxn_opcodes_h_l2265_c7_2b90
n8_MUX_uxn_opcodes_h_l2265_c7_2b90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2265_c7_2b90_cond,
n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue,
n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse,
n8_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output);

-- t16_MUX_uxn_opcodes_h_l2265_c7_2b90
t16_MUX_uxn_opcodes_h_l2265_c7_2b90 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2265_c7_2b90_cond,
t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue,
t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse,
t16_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90
result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond,
result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90
result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond,
result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90
result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90
result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90
result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11
BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_left,
BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_right,
BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output);

-- n8_MUX_uxn_opcodes_h_l2268_c7_fe9f
n8_MUX_uxn_opcodes_h_l2268_c7_fe9f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond,
n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue,
n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse,
n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output);

-- t16_MUX_uxn_opcodes_h_l2268_c7_fe9f
t16_MUX_uxn_opcodes_h_l2268_c7_fe9f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond,
t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue,
t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse,
t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f
result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond,
result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f
result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f
result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f
result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2270_c3_051f
CONST_SL_8_uxn_opcodes_h_l2270_c3_051f : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_x,
CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429
BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_left,
BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_right,
BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output);

-- n8_MUX_uxn_opcodes_h_l2273_c7_1ce9
n8_MUX_uxn_opcodes_h_l2273_c7_1ce9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond,
n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue,
n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse,
n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output);

-- t16_MUX_uxn_opcodes_h_l2273_c7_1ce9
t16_MUX_uxn_opcodes_h_l2273_c7_1ce9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond,
t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue,
t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse,
t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9
result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond,
result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9
result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9
result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9
result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee
BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_left,
BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_right,
BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1
BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_left,
BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_right,
BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output);

-- n8_MUX_uxn_opcodes_h_l2276_c7_531c
n8_MUX_uxn_opcodes_h_l2276_c7_531c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2276_c7_531c_cond,
n8_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue,
n8_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse,
n8_MUX_uxn_opcodes_h_l2276_c7_531c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c
result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond,
result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c
result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c
result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c
result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2279_c30_c336
sp_relative_shift_uxn_opcodes_h_l2279_c30_c336 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_ins,
sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_x,
sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_y,
sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771
BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_left,
BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_right,
BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f
result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f
result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output,
 n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
 t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output,
 n8_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output,
 t16_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output,
 n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output,
 t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output,
 CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output,
 n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output,
 t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output,
 n8_MUX_uxn_opcodes_h_l2276_c7_531c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2262_c3_2a1e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2266_c3_6e7f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2271_c3_b727 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2268_c7_fe9f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2285_c3_28c3 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_94be_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_d85a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_5206_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_a9ce_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2284_l2276_l2273_l2268_l2265_DUPLICATE_4d69_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2274_l2269_DUPLICATE_cd25_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_7ccb_uxn_opcodes_h_l2290_l2253_DUPLICATE_60d9_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2266_c3_6e7f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2266_c3_6e7f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2271_c3_b727 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2271_c3_b727;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_right := to_unsigned(4, 3);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_y := resize(to_signed(-3, 3), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2262_c3_2a1e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2262_c3_2a1e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2285_c3_28c3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2285_c3_28c3;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l2276_c11_43e1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2274_l2269_DUPLICATE_cd25 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2274_l2269_DUPLICATE_cd25_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2284_l2276_l2273_l2268_l2265_DUPLICATE_4d69 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2284_l2276_l2273_l2268_l2265_DUPLICATE_4d69_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_a9ce LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_a9ce_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2265_c11_d60e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2273_c11_2429] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_left;
     BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output := BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2279_c30_c336] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_ins;
     sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_x;
     sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_return_output := sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2284_c11_d771] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_left;
     BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output := BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_d85a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_d85a_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_5206 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_5206_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2258_c6_d2c6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2268_c11_cb11] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_left;
     BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output := BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2268_c7_fe9f_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_94be LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_94be_return_output := result.u16_value;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2258_c6_d2c6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2265_c11_d60e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2268_c11_cb11_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2273_c11_2429_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2276_c11_43e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2284_c11_d771_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2274_l2269_DUPLICATE_cd25_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2274_l2269_DUPLICATE_cd25_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_5206_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_5206_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_5206_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_5206_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_5206_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_94be_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_94be_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_94be_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_94be_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_94be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2284_l2276_l2273_l2268_l2265_DUPLICATE_4d69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2284_l2276_l2273_l2268_l2265_DUPLICATE_4d69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2284_l2276_l2273_l2268_l2265_DUPLICATE_4d69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2284_l2276_l2273_l2268_l2265_DUPLICATE_4d69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2284_l2276_l2273_l2268_l2265_DUPLICATE_4d69_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_a9ce_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_a9ce_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_a9ce_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_a9ce_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2284_l2273_l2268_l2265_l2258_DUPLICATE_a9ce_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_d85a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_d85a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_d85a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_d85a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2276_l2273_l2268_l2265_l2258_DUPLICATE_d85a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2279_c30_c336_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2284_c7_ea4f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2270_c3_051f] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_return_output := CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2274_c3_b7ee] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_left;
     BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_return_output := BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2276_c7_531c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2284_c7_ea4f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2276_c7_531c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output := result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2284_c7_ea4f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2276_c7_531c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2276_c7_531c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_cond;
     n8_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue;
     n8_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_return_output := n8_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2274_c3_b7ee_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2270_c3_051f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2284_c7_ea4f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2273_c7_1ce9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output := result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2273_c7_1ce9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2265_c7_2b90] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2276_c7_531c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;

     -- t16_MUX[uxn_opcodes_h_l2273_c7_1ce9] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond <= VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond;
     t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue;
     t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output := t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2276_c7_531c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2273_c7_1ce9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond;
     n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue;
     n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output := n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2276_c7_531c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2276_c7_531c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2273_c7_1ce9] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2273_c7_1ce9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond;
     n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue;
     n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output := n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;

     -- t16_MUX[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond <= VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond;
     t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue;
     t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output := t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2258_c2_8d8f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2273_c7_1ce9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output := result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2273_c7_1ce9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2265_c7_2b90] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output := result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;

     -- t16_MUX[uxn_opcodes_h_l2265_c7_2b90] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2265_c7_2b90_cond <= VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_cond;
     t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue;
     t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output := t16_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;

     -- n8_MUX[uxn_opcodes_h_l2265_c7_2b90] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2265_c7_2b90_cond <= VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_cond;
     n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue;
     n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output := n8_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2265_c7_2b90] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output := result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2268_c7_fe9f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2268_c7_fe9f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l2265_c7_2b90] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;

     -- t16_MUX[uxn_opcodes_h_l2258_c2_8d8f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond <= VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond;
     t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue;
     t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output := t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2258_c2_8d8f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output := result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2258_c2_8d8f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2258_c2_8d8f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond;
     n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue;
     n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output := n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2265_c7_2b90] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2265_c7_2b90] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2265_c7_2b90_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2258_c2_8d8f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2258_c2_8d8f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2258_c2_8d8f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_7ccb_uxn_opcodes_h_l2290_l2253_DUPLICATE_60d9 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_7ccb_uxn_opcodes_h_l2290_l2253_DUPLICATE_60d9_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_7ccb(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2258_c2_8d8f_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_7ccb_uxn_opcodes_h_l2290_l2253_DUPLICATE_60d9_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_7ccb_uxn_opcodes_h_l2290_l2253_DUPLICATE_60d9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
