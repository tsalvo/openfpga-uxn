-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity eor2_0CLK_06b39b76 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end eor2_0CLK_06b39b76;
architecture arch of eor2_0CLK_06b39b76 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1023_c6_3b71]
signal BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1023_c2_2188]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1023_c2_2188]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1023_c2_2188]
signal result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1023_c2_2188]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1023_c2_2188]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1023_c2_2188]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1023_c2_2188]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1023_c2_2188]
signal n16_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1023_c2_2188]
signal tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1023_c2_2188]
signal t16_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1031_c11_e268]
signal BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1031_c7_97df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1031_c7_97df]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1031_c7_97df]
signal result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1031_c7_97df]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1031_c7_97df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1031_c7_97df]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1031_c7_97df]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1031_c7_97df]
signal n16_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1031_c7_97df]
signal tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1031_c7_97df]
signal t16_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1034_c11_516a]
signal BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1034_c7_c2b9]
signal t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1037_c30_a8c2]
signal sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1039_c11_ddba]
signal BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1039_c7_abc3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1039_c7_abc3]
signal result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1039_c7_abc3]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1039_c7_abc3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1039_c7_abc3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1039_c7_abc3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l1039_c7_abc3]
signal n16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(15 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l1039_c7_abc3]
signal tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(15 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1041_c11_3f5f]
signal BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_left : unsigned(15 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_right : unsigned(15 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1047_c11_1730]
signal BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1047_c7_17ea]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1047_c7_17ea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1047_c7_17ea]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71
BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_left,
BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_right,
BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188
result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188
result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- n16_MUX_uxn_opcodes_h_l1023_c2_2188
n16_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
n16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
n16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
n16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1023_c2_2188
tmp16_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- t16_MUX_uxn_opcodes_h_l1023_c2_2188
t16_MUX_uxn_opcodes_h_l1023_c2_2188 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1023_c2_2188_cond,
t16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue,
t16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse,
t16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268
BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_left,
BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_right,
BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df
result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df
result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df
result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df
result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df
result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- n16_MUX_uxn_opcodes_h_l1031_c7_97df
n16_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
n16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
n16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
n16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1031_c7_97df
tmp16_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- t16_MUX_uxn_opcodes_h_l1031_c7_97df
t16_MUX_uxn_opcodes_h_l1031_c7_97df : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1031_c7_97df_cond,
t16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue,
t16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse,
t16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a
BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_left,
BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_right,
BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9
result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9
result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9
result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9
result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- n16_MUX_uxn_opcodes_h_l1034_c7_c2b9
n16_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9
tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- t16_MUX_uxn_opcodes_h_l1034_c7_c2b9
t16_MUX_uxn_opcodes_h_l1034_c7_c2b9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond,
t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue,
t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse,
t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2
sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_ins,
sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_x,
sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_y,
sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba
BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_left,
BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_right,
BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3
result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_cond,
result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output);

-- n16_MUX_uxn_opcodes_h_l1039_c7_abc3
n16_MUX_uxn_opcodes_h_l1039_c7_abc3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond,
n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue,
n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse,
n16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output);

-- tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3
tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond,
tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue,
tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse,
tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f
BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f : entity work.BIN_OP_XOR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_left,
BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_right,
BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730
BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_left,
BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_right,
BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea
result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea
result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 n16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 t16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 n16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 t16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output,
 sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output,
 n16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output,
 tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1028_c3_bebb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1032_c3_35d4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1044_c3_27bc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1023_l1039_l1031_DUPLICATE_0eda_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1034_l1023_l1039_l1031_DUPLICATE_0a50_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1034_l1023_l1031_DUPLICATE_20ed_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1034_l1023_l1031_l1047_DUPLICATE_bd2a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_0909_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_a0ad_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1034_l1039_DUPLICATE_0877_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1053_l1019_DUPLICATE_58f2_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1028_c3_bebb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1028_c3_bebb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_right := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1032_c3_35d4 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1032_c3_35d4;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1044_c3_27bc := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1044_c3_27bc;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := t16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l1047_c11_1730] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_left;
     BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output := BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1023_c6_3b71] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_left;
     BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output := BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_0909 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_0909_return_output := result.is_stack_operation_16bit;

     -- sp_relative_shift[uxn_opcodes_h_l1037_c30_a8c2] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_ins;
     sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_x;
     sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_return_output := sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1034_l1023_l1031_DUPLICATE_20ed LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1034_l1023_l1031_DUPLICATE_20ed_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1031_c11_e268] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_left;
     BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output := BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_a0ad LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_a0ad_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1034_l1039_DUPLICATE_0877 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1034_l1039_DUPLICATE_0877_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1034_l1023_l1031_l1047_DUPLICATE_bd2a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1034_l1023_l1031_l1047_DUPLICATE_bd2a_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1034_c11_516a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1039_c11_ddba] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_left;
     BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output := BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;

     -- BIN_OP_XOR[uxn_opcodes_h_l1041_c11_3f5f] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_left;
     BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_return_output := BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1023_l1039_l1031_DUPLICATE_0eda LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1023_l1039_l1031_DUPLICATE_0eda_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1034_l1023_l1039_l1031_DUPLICATE_0a50 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1034_l1023_l1039_l1031_DUPLICATE_0a50_return_output := result.u16_value;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1023_c6_3b71_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1031_c11_e268_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1034_c11_516a_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1039_c11_ddba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1047_c11_1730_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1041_c11_3f5f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1034_l1023_l1031_DUPLICATE_20ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1034_l1023_l1031_DUPLICATE_20ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1034_l1023_l1031_DUPLICATE_20ed_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1034_l1023_l1039_l1031_DUPLICATE_0a50_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1034_l1023_l1039_l1031_DUPLICATE_0a50_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1034_l1023_l1039_l1031_DUPLICATE_0a50_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1034_l1023_l1039_l1031_DUPLICATE_0a50_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_a0ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_a0ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_a0ad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_a0ad_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1023_l1039_l1031_DUPLICATE_0eda_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1023_l1039_l1031_DUPLICATE_0eda_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1023_l1039_l1031_DUPLICATE_0eda_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_0909_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_0909_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_0909_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1034_l1039_l1031_l1047_DUPLICATE_0909_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1034_l1023_l1031_l1047_DUPLICATE_bd2a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1034_l1023_l1031_l1047_DUPLICATE_bd2a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1034_l1023_l1031_l1047_DUPLICATE_bd2a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1034_l1023_l1031_l1047_DUPLICATE_bd2a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1034_l1039_DUPLICATE_0877_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1034_l1039_DUPLICATE_0877_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1037_c30_a8c2_return_output;
     -- t16_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1039_c7_abc3] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond;
     tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output := tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;

     -- n16_MUX[uxn_opcodes_h_l1039_c7_abc3] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond <= VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_cond;
     n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue;
     n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output := n16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1039_c7_abc3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output := result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1039_c7_abc3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1039_c7_abc3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1047_c7_17ea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1047_c7_17ea] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1047_c7_17ea] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- Submodule level 2
     VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1047_c7_17ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1039_c7_abc3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- n16_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1039_c7_abc3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1039_c7_abc3] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- t16_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     t16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     t16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := t16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1039_c7_abc3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     -- t16_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     t16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     t16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := t16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- n16_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     n16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     n16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := n16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1034_c7_c2b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1034_c7_c2b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- n16_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     n16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     n16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := n16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1031_c7_97df] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1031_c7_97df_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1023_c2_2188] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1053_l1019_DUPLICATE_58f2 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1053_l1019_DUPLICATE_58f2_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1023_c2_2188_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1023_c2_2188_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1053_l1019_DUPLICATE_58f2_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l1053_l1019_DUPLICATE_58f2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
