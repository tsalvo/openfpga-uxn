-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 134
entity uint8_mux128_0CLK_9347d63d is
port(
 sel : in unsigned(6 downto 0);
 in0 : in unsigned(7 downto 0);
 in1 : in unsigned(7 downto 0);
 in2 : in unsigned(7 downto 0);
 in3 : in unsigned(7 downto 0);
 in4 : in unsigned(7 downto 0);
 in5 : in unsigned(7 downto 0);
 in6 : in unsigned(7 downto 0);
 in7 : in unsigned(7 downto 0);
 in8 : in unsigned(7 downto 0);
 in9 : in unsigned(7 downto 0);
 in10 : in unsigned(7 downto 0);
 in11 : in unsigned(7 downto 0);
 in12 : in unsigned(7 downto 0);
 in13 : in unsigned(7 downto 0);
 in14 : in unsigned(7 downto 0);
 in15 : in unsigned(7 downto 0);
 in16 : in unsigned(7 downto 0);
 in17 : in unsigned(7 downto 0);
 in18 : in unsigned(7 downto 0);
 in19 : in unsigned(7 downto 0);
 in20 : in unsigned(7 downto 0);
 in21 : in unsigned(7 downto 0);
 in22 : in unsigned(7 downto 0);
 in23 : in unsigned(7 downto 0);
 in24 : in unsigned(7 downto 0);
 in25 : in unsigned(7 downto 0);
 in26 : in unsigned(7 downto 0);
 in27 : in unsigned(7 downto 0);
 in28 : in unsigned(7 downto 0);
 in29 : in unsigned(7 downto 0);
 in30 : in unsigned(7 downto 0);
 in31 : in unsigned(7 downto 0);
 in32 : in unsigned(7 downto 0);
 in33 : in unsigned(7 downto 0);
 in34 : in unsigned(7 downto 0);
 in35 : in unsigned(7 downto 0);
 in36 : in unsigned(7 downto 0);
 in37 : in unsigned(7 downto 0);
 in38 : in unsigned(7 downto 0);
 in39 : in unsigned(7 downto 0);
 in40 : in unsigned(7 downto 0);
 in41 : in unsigned(7 downto 0);
 in42 : in unsigned(7 downto 0);
 in43 : in unsigned(7 downto 0);
 in44 : in unsigned(7 downto 0);
 in45 : in unsigned(7 downto 0);
 in46 : in unsigned(7 downto 0);
 in47 : in unsigned(7 downto 0);
 in48 : in unsigned(7 downto 0);
 in49 : in unsigned(7 downto 0);
 in50 : in unsigned(7 downto 0);
 in51 : in unsigned(7 downto 0);
 in52 : in unsigned(7 downto 0);
 in53 : in unsigned(7 downto 0);
 in54 : in unsigned(7 downto 0);
 in55 : in unsigned(7 downto 0);
 in56 : in unsigned(7 downto 0);
 in57 : in unsigned(7 downto 0);
 in58 : in unsigned(7 downto 0);
 in59 : in unsigned(7 downto 0);
 in60 : in unsigned(7 downto 0);
 in61 : in unsigned(7 downto 0);
 in62 : in unsigned(7 downto 0);
 in63 : in unsigned(7 downto 0);
 in64 : in unsigned(7 downto 0);
 in65 : in unsigned(7 downto 0);
 in66 : in unsigned(7 downto 0);
 in67 : in unsigned(7 downto 0);
 in68 : in unsigned(7 downto 0);
 in69 : in unsigned(7 downto 0);
 in70 : in unsigned(7 downto 0);
 in71 : in unsigned(7 downto 0);
 in72 : in unsigned(7 downto 0);
 in73 : in unsigned(7 downto 0);
 in74 : in unsigned(7 downto 0);
 in75 : in unsigned(7 downto 0);
 in76 : in unsigned(7 downto 0);
 in77 : in unsigned(7 downto 0);
 in78 : in unsigned(7 downto 0);
 in79 : in unsigned(7 downto 0);
 in80 : in unsigned(7 downto 0);
 in81 : in unsigned(7 downto 0);
 in82 : in unsigned(7 downto 0);
 in83 : in unsigned(7 downto 0);
 in84 : in unsigned(7 downto 0);
 in85 : in unsigned(7 downto 0);
 in86 : in unsigned(7 downto 0);
 in87 : in unsigned(7 downto 0);
 in88 : in unsigned(7 downto 0);
 in89 : in unsigned(7 downto 0);
 in90 : in unsigned(7 downto 0);
 in91 : in unsigned(7 downto 0);
 in92 : in unsigned(7 downto 0);
 in93 : in unsigned(7 downto 0);
 in94 : in unsigned(7 downto 0);
 in95 : in unsigned(7 downto 0);
 in96 : in unsigned(7 downto 0);
 in97 : in unsigned(7 downto 0);
 in98 : in unsigned(7 downto 0);
 in99 : in unsigned(7 downto 0);
 in100 : in unsigned(7 downto 0);
 in101 : in unsigned(7 downto 0);
 in102 : in unsigned(7 downto 0);
 in103 : in unsigned(7 downto 0);
 in104 : in unsigned(7 downto 0);
 in105 : in unsigned(7 downto 0);
 in106 : in unsigned(7 downto 0);
 in107 : in unsigned(7 downto 0);
 in108 : in unsigned(7 downto 0);
 in109 : in unsigned(7 downto 0);
 in110 : in unsigned(7 downto 0);
 in111 : in unsigned(7 downto 0);
 in112 : in unsigned(7 downto 0);
 in113 : in unsigned(7 downto 0);
 in114 : in unsigned(7 downto 0);
 in115 : in unsigned(7 downto 0);
 in116 : in unsigned(7 downto 0);
 in117 : in unsigned(7 downto 0);
 in118 : in unsigned(7 downto 0);
 in119 : in unsigned(7 downto 0);
 in120 : in unsigned(7 downto 0);
 in121 : in unsigned(7 downto 0);
 in122 : in unsigned(7 downto 0);
 in123 : in unsigned(7 downto 0);
 in124 : in unsigned(7 downto 0);
 in125 : in unsigned(7 downto 0);
 in126 : in unsigned(7 downto 0);
 in127 : in unsigned(7 downto 0);
 return_output : out unsigned(7 downto 0));
end uint8_mux128_0CLK_9347d63d;
architecture arch of uint8_mux128_0CLK_9347d63d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_70c7]
signal layer0_node0_MUX_bit_math_h_l18_c3_70c7_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_70c7_iftrue : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_70c7_iffalse : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_70c7_return_output : unsigned(7 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_dc12]
signal layer0_node1_MUX_bit_math_h_l29_c3_dc12_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_dc12_iftrue : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_dc12_iffalse : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_dc12_return_output : unsigned(7 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_3404]
signal layer0_node2_MUX_bit_math_h_l40_c3_3404_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_3404_iftrue : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_3404_iffalse : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_3404_return_output : unsigned(7 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_cc01]
signal layer0_node3_MUX_bit_math_h_l51_c3_cc01_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_cc01_iftrue : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_cc01_iffalse : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_cc01_return_output : unsigned(7 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_7793]
signal layer0_node4_MUX_bit_math_h_l62_c3_7793_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_7793_iftrue : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_7793_iffalse : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_7793_return_output : unsigned(7 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_2acd]
signal layer0_node5_MUX_bit_math_h_l73_c3_2acd_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_2acd_iftrue : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_2acd_iffalse : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_2acd_return_output : unsigned(7 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_494b]
signal layer0_node6_MUX_bit_math_h_l84_c3_494b_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_494b_iftrue : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_494b_iffalse : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_494b_return_output : unsigned(7 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_daab]
signal layer0_node7_MUX_bit_math_h_l95_c3_daab_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_daab_iftrue : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_daab_iffalse : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_daab_return_output : unsigned(7 downto 0);

-- layer0_node8_MUX[bit_math_h_l106_c3_d50d]
signal layer0_node8_MUX_bit_math_h_l106_c3_d50d_cond : unsigned(0 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_d50d_iftrue : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_d50d_iffalse : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_d50d_return_output : unsigned(7 downto 0);

-- layer0_node9_MUX[bit_math_h_l117_c3_c9ee]
signal layer0_node9_MUX_bit_math_h_l117_c3_c9ee_cond : unsigned(0 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iftrue : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iffalse : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_c9ee_return_output : unsigned(7 downto 0);

-- layer0_node10_MUX[bit_math_h_l128_c3_06d1]
signal layer0_node10_MUX_bit_math_h_l128_c3_06d1_cond : unsigned(0 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_06d1_iftrue : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_06d1_iffalse : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_06d1_return_output : unsigned(7 downto 0);

-- layer0_node11_MUX[bit_math_h_l139_c3_13dc]
signal layer0_node11_MUX_bit_math_h_l139_c3_13dc_cond : unsigned(0 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_13dc_iftrue : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_13dc_iffalse : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_13dc_return_output : unsigned(7 downto 0);

-- layer0_node12_MUX[bit_math_h_l150_c3_af2c]
signal layer0_node12_MUX_bit_math_h_l150_c3_af2c_cond : unsigned(0 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_af2c_iftrue : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_af2c_iffalse : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_af2c_return_output : unsigned(7 downto 0);

-- layer0_node13_MUX[bit_math_h_l161_c3_c865]
signal layer0_node13_MUX_bit_math_h_l161_c3_c865_cond : unsigned(0 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_c865_iftrue : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_c865_iffalse : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_c865_return_output : unsigned(7 downto 0);

-- layer0_node14_MUX[bit_math_h_l172_c3_1937]
signal layer0_node14_MUX_bit_math_h_l172_c3_1937_cond : unsigned(0 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_1937_iftrue : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_1937_iffalse : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_1937_return_output : unsigned(7 downto 0);

-- layer0_node15_MUX[bit_math_h_l183_c3_6211]
signal layer0_node15_MUX_bit_math_h_l183_c3_6211_cond : unsigned(0 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_6211_iftrue : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_6211_iffalse : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_6211_return_output : unsigned(7 downto 0);

-- layer0_node16_MUX[bit_math_h_l194_c3_6e24]
signal layer0_node16_MUX_bit_math_h_l194_c3_6e24_cond : unsigned(0 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_6e24_iftrue : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_6e24_iffalse : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_6e24_return_output : unsigned(7 downto 0);

-- layer0_node17_MUX[bit_math_h_l205_c3_4b2c]
signal layer0_node17_MUX_bit_math_h_l205_c3_4b2c_cond : unsigned(0 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iftrue : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iffalse : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_4b2c_return_output : unsigned(7 downto 0);

-- layer0_node18_MUX[bit_math_h_l216_c3_0b83]
signal layer0_node18_MUX_bit_math_h_l216_c3_0b83_cond : unsigned(0 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_0b83_iftrue : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_0b83_iffalse : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_0b83_return_output : unsigned(7 downto 0);

-- layer0_node19_MUX[bit_math_h_l227_c3_1e36]
signal layer0_node19_MUX_bit_math_h_l227_c3_1e36_cond : unsigned(0 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1e36_iftrue : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1e36_iffalse : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_1e36_return_output : unsigned(7 downto 0);

-- layer0_node20_MUX[bit_math_h_l238_c3_5458]
signal layer0_node20_MUX_bit_math_h_l238_c3_5458_cond : unsigned(0 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_5458_iftrue : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_5458_iffalse : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_5458_return_output : unsigned(7 downto 0);

-- layer0_node21_MUX[bit_math_h_l249_c3_c173]
signal layer0_node21_MUX_bit_math_h_l249_c3_c173_cond : unsigned(0 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_c173_iftrue : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_c173_iffalse : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_c173_return_output : unsigned(7 downto 0);

-- layer0_node22_MUX[bit_math_h_l260_c3_fce5]
signal layer0_node22_MUX_bit_math_h_l260_c3_fce5_cond : unsigned(0 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_fce5_iftrue : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_fce5_iffalse : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_fce5_return_output : unsigned(7 downto 0);

-- layer0_node23_MUX[bit_math_h_l271_c3_a82d]
signal layer0_node23_MUX_bit_math_h_l271_c3_a82d_cond : unsigned(0 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_a82d_iftrue : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_a82d_iffalse : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_a82d_return_output : unsigned(7 downto 0);

-- layer0_node24_MUX[bit_math_h_l282_c3_6611]
signal layer0_node24_MUX_bit_math_h_l282_c3_6611_cond : unsigned(0 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_6611_iftrue : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_6611_iffalse : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_6611_return_output : unsigned(7 downto 0);

-- layer0_node25_MUX[bit_math_h_l293_c3_b4b9]
signal layer0_node25_MUX_bit_math_h_l293_c3_b4b9_cond : unsigned(0 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iftrue : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iffalse : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_b4b9_return_output : unsigned(7 downto 0);

-- layer0_node26_MUX[bit_math_h_l304_c3_2bce]
signal layer0_node26_MUX_bit_math_h_l304_c3_2bce_cond : unsigned(0 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_2bce_iftrue : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_2bce_iffalse : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_2bce_return_output : unsigned(7 downto 0);

-- layer0_node27_MUX[bit_math_h_l315_c3_7789]
signal layer0_node27_MUX_bit_math_h_l315_c3_7789_cond : unsigned(0 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_7789_iftrue : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_7789_iffalse : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_7789_return_output : unsigned(7 downto 0);

-- layer0_node28_MUX[bit_math_h_l326_c3_098d]
signal layer0_node28_MUX_bit_math_h_l326_c3_098d_cond : unsigned(0 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_098d_iftrue : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_098d_iffalse : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_098d_return_output : unsigned(7 downto 0);

-- layer0_node29_MUX[bit_math_h_l337_c3_9c87]
signal layer0_node29_MUX_bit_math_h_l337_c3_9c87_cond : unsigned(0 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_9c87_iftrue : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_9c87_iffalse : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_9c87_return_output : unsigned(7 downto 0);

-- layer0_node30_MUX[bit_math_h_l348_c3_6b0d]
signal layer0_node30_MUX_bit_math_h_l348_c3_6b0d_cond : unsigned(0 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iftrue : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iffalse : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_6b0d_return_output : unsigned(7 downto 0);

-- layer0_node31_MUX[bit_math_h_l359_c3_5065]
signal layer0_node31_MUX_bit_math_h_l359_c3_5065_cond : unsigned(0 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_5065_iftrue : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_5065_iffalse : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_5065_return_output : unsigned(7 downto 0);

-- layer0_node32_MUX[bit_math_h_l370_c3_4893]
signal layer0_node32_MUX_bit_math_h_l370_c3_4893_cond : unsigned(0 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_4893_iftrue : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_4893_iffalse : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_4893_return_output : unsigned(7 downto 0);

-- layer0_node33_MUX[bit_math_h_l381_c3_8132]
signal layer0_node33_MUX_bit_math_h_l381_c3_8132_cond : unsigned(0 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_8132_iftrue : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_8132_iffalse : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_8132_return_output : unsigned(7 downto 0);

-- layer0_node34_MUX[bit_math_h_l392_c3_59bd]
signal layer0_node34_MUX_bit_math_h_l392_c3_59bd_cond : unsigned(0 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_59bd_iftrue : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_59bd_iffalse : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_59bd_return_output : unsigned(7 downto 0);

-- layer0_node35_MUX[bit_math_h_l403_c3_6326]
signal layer0_node35_MUX_bit_math_h_l403_c3_6326_cond : unsigned(0 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_6326_iftrue : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_6326_iffalse : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_6326_return_output : unsigned(7 downto 0);

-- layer0_node36_MUX[bit_math_h_l414_c3_7348]
signal layer0_node36_MUX_bit_math_h_l414_c3_7348_cond : unsigned(0 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_7348_iftrue : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_7348_iffalse : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_7348_return_output : unsigned(7 downto 0);

-- layer0_node37_MUX[bit_math_h_l425_c3_f929]
signal layer0_node37_MUX_bit_math_h_l425_c3_f929_cond : unsigned(0 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_f929_iftrue : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_f929_iffalse : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_f929_return_output : unsigned(7 downto 0);

-- layer0_node38_MUX[bit_math_h_l436_c3_d3a0]
signal layer0_node38_MUX_bit_math_h_l436_c3_d3a0_cond : unsigned(0 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iftrue : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iffalse : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_d3a0_return_output : unsigned(7 downto 0);

-- layer0_node39_MUX[bit_math_h_l447_c3_7b35]
signal layer0_node39_MUX_bit_math_h_l447_c3_7b35_cond : unsigned(0 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_7b35_iftrue : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_7b35_iffalse : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_7b35_return_output : unsigned(7 downto 0);

-- layer0_node40_MUX[bit_math_h_l458_c3_426b]
signal layer0_node40_MUX_bit_math_h_l458_c3_426b_cond : unsigned(0 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_426b_iftrue : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_426b_iffalse : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_426b_return_output : unsigned(7 downto 0);

-- layer0_node41_MUX[bit_math_h_l469_c3_47d5]
signal layer0_node41_MUX_bit_math_h_l469_c3_47d5_cond : unsigned(0 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_47d5_iftrue : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_47d5_iffalse : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_47d5_return_output : unsigned(7 downto 0);

-- layer0_node42_MUX[bit_math_h_l480_c3_50c3]
signal layer0_node42_MUX_bit_math_h_l480_c3_50c3_cond : unsigned(0 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_50c3_iftrue : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_50c3_iffalse : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_50c3_return_output : unsigned(7 downto 0);

-- layer0_node43_MUX[bit_math_h_l491_c3_6ed7]
signal layer0_node43_MUX_bit_math_h_l491_c3_6ed7_cond : unsigned(0 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iftrue : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iffalse : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_6ed7_return_output : unsigned(7 downto 0);

-- layer0_node44_MUX[bit_math_h_l502_c3_84a4]
signal layer0_node44_MUX_bit_math_h_l502_c3_84a4_cond : unsigned(0 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_84a4_iftrue : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_84a4_iffalse : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_84a4_return_output : unsigned(7 downto 0);

-- layer0_node45_MUX[bit_math_h_l513_c3_552e]
signal layer0_node45_MUX_bit_math_h_l513_c3_552e_cond : unsigned(0 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_552e_iftrue : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_552e_iffalse : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_552e_return_output : unsigned(7 downto 0);

-- layer0_node46_MUX[bit_math_h_l524_c3_42cd]
signal layer0_node46_MUX_bit_math_h_l524_c3_42cd_cond : unsigned(0 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_42cd_iftrue : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_42cd_iffalse : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_42cd_return_output : unsigned(7 downto 0);

-- layer0_node47_MUX[bit_math_h_l535_c3_18b2]
signal layer0_node47_MUX_bit_math_h_l535_c3_18b2_cond : unsigned(0 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_18b2_iftrue : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_18b2_iffalse : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_18b2_return_output : unsigned(7 downto 0);

-- layer0_node48_MUX[bit_math_h_l546_c3_e9fe]
signal layer0_node48_MUX_bit_math_h_l546_c3_e9fe_cond : unsigned(0 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iftrue : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iffalse : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_e9fe_return_output : unsigned(7 downto 0);

-- layer0_node49_MUX[bit_math_h_l557_c3_68c1]
signal layer0_node49_MUX_bit_math_h_l557_c3_68c1_cond : unsigned(0 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_68c1_iftrue : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_68c1_iffalse : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_68c1_return_output : unsigned(7 downto 0);

-- layer0_node50_MUX[bit_math_h_l568_c3_8ec7]
signal layer0_node50_MUX_bit_math_h_l568_c3_8ec7_cond : unsigned(0 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iftrue : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iffalse : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_8ec7_return_output : unsigned(7 downto 0);

-- layer0_node51_MUX[bit_math_h_l579_c3_5985]
signal layer0_node51_MUX_bit_math_h_l579_c3_5985_cond : unsigned(0 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_5985_iftrue : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_5985_iffalse : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_5985_return_output : unsigned(7 downto 0);

-- layer0_node52_MUX[bit_math_h_l590_c3_90c2]
signal layer0_node52_MUX_bit_math_h_l590_c3_90c2_cond : unsigned(0 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_90c2_iftrue : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_90c2_iffalse : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_90c2_return_output : unsigned(7 downto 0);

-- layer0_node53_MUX[bit_math_h_l601_c3_5a9e]
signal layer0_node53_MUX_bit_math_h_l601_c3_5a9e_cond : unsigned(0 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iftrue : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iffalse : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_5a9e_return_output : unsigned(7 downto 0);

-- layer0_node54_MUX[bit_math_h_l612_c3_235a]
signal layer0_node54_MUX_bit_math_h_l612_c3_235a_cond : unsigned(0 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_235a_iftrue : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_235a_iffalse : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_235a_return_output : unsigned(7 downto 0);

-- layer0_node55_MUX[bit_math_h_l623_c3_1dea]
signal layer0_node55_MUX_bit_math_h_l623_c3_1dea_cond : unsigned(0 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_1dea_iftrue : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_1dea_iffalse : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_1dea_return_output : unsigned(7 downto 0);

-- layer0_node56_MUX[bit_math_h_l634_c3_f6e3]
signal layer0_node56_MUX_bit_math_h_l634_c3_f6e3_cond : unsigned(0 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iftrue : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iffalse : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_f6e3_return_output : unsigned(7 downto 0);

-- layer0_node57_MUX[bit_math_h_l645_c3_eeb0]
signal layer0_node57_MUX_bit_math_h_l645_c3_eeb0_cond : unsigned(0 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iftrue : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iffalse : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_eeb0_return_output : unsigned(7 downto 0);

-- layer0_node58_MUX[bit_math_h_l656_c3_b995]
signal layer0_node58_MUX_bit_math_h_l656_c3_b995_cond : unsigned(0 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_b995_iftrue : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_b995_iffalse : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_b995_return_output : unsigned(7 downto 0);

-- layer0_node59_MUX[bit_math_h_l667_c3_b104]
signal layer0_node59_MUX_bit_math_h_l667_c3_b104_cond : unsigned(0 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_b104_iftrue : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_b104_iffalse : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_b104_return_output : unsigned(7 downto 0);

-- layer0_node60_MUX[bit_math_h_l678_c3_7571]
signal layer0_node60_MUX_bit_math_h_l678_c3_7571_cond : unsigned(0 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_7571_iftrue : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_7571_iffalse : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_7571_return_output : unsigned(7 downto 0);

-- layer0_node61_MUX[bit_math_h_l689_c3_580e]
signal layer0_node61_MUX_bit_math_h_l689_c3_580e_cond : unsigned(0 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_580e_iftrue : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_580e_iffalse : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_580e_return_output : unsigned(7 downto 0);

-- layer0_node62_MUX[bit_math_h_l700_c3_9f5f]
signal layer0_node62_MUX_bit_math_h_l700_c3_9f5f_cond : unsigned(0 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iftrue : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iffalse : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_9f5f_return_output : unsigned(7 downto 0);

-- layer0_node63_MUX[bit_math_h_l711_c3_17f2]
signal layer0_node63_MUX_bit_math_h_l711_c3_17f2_cond : unsigned(0 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_17f2_iftrue : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_17f2_iffalse : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_17f2_return_output : unsigned(7 downto 0);

-- layer1_node0_MUX[bit_math_h_l728_c3_23e3]
signal layer1_node0_MUX_bit_math_h_l728_c3_23e3_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_23e3_iftrue : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_23e3_iffalse : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_23e3_return_output : unsigned(7 downto 0);

-- layer1_node1_MUX[bit_math_h_l739_c3_57f6]
signal layer1_node1_MUX_bit_math_h_l739_c3_57f6_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_57f6_iftrue : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_57f6_iffalse : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_57f6_return_output : unsigned(7 downto 0);

-- layer1_node2_MUX[bit_math_h_l750_c3_b86b]
signal layer1_node2_MUX_bit_math_h_l750_c3_b86b_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_b86b_iftrue : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_b86b_iffalse : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_b86b_return_output : unsigned(7 downto 0);

-- layer1_node3_MUX[bit_math_h_l761_c3_2586]
signal layer1_node3_MUX_bit_math_h_l761_c3_2586_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_2586_iftrue : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_2586_iffalse : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_2586_return_output : unsigned(7 downto 0);

-- layer1_node4_MUX[bit_math_h_l772_c3_857f]
signal layer1_node4_MUX_bit_math_h_l772_c3_857f_cond : unsigned(0 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_857f_iftrue : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_857f_iffalse : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_857f_return_output : unsigned(7 downto 0);

-- layer1_node5_MUX[bit_math_h_l783_c3_f8bc]
signal layer1_node5_MUX_bit_math_h_l783_c3_f8bc_cond : unsigned(0 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iftrue : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iffalse : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_f8bc_return_output : unsigned(7 downto 0);

-- layer1_node6_MUX[bit_math_h_l794_c3_f4dd]
signal layer1_node6_MUX_bit_math_h_l794_c3_f4dd_cond : unsigned(0 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iftrue : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iffalse : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_f4dd_return_output : unsigned(7 downto 0);

-- layer1_node7_MUX[bit_math_h_l805_c3_e535]
signal layer1_node7_MUX_bit_math_h_l805_c3_e535_cond : unsigned(0 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_e535_iftrue : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_e535_iffalse : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_e535_return_output : unsigned(7 downto 0);

-- layer1_node8_MUX[bit_math_h_l816_c3_e51d]
signal layer1_node8_MUX_bit_math_h_l816_c3_e51d_cond : unsigned(0 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_e51d_iftrue : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_e51d_iffalse : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_e51d_return_output : unsigned(7 downto 0);

-- layer1_node9_MUX[bit_math_h_l827_c3_4f17]
signal layer1_node9_MUX_bit_math_h_l827_c3_4f17_cond : unsigned(0 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_4f17_iftrue : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_4f17_iffalse : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_4f17_return_output : unsigned(7 downto 0);

-- layer1_node10_MUX[bit_math_h_l838_c3_8caa]
signal layer1_node10_MUX_bit_math_h_l838_c3_8caa_cond : unsigned(0 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_8caa_iftrue : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_8caa_iffalse : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_8caa_return_output : unsigned(7 downto 0);

-- layer1_node11_MUX[bit_math_h_l849_c3_c418]
signal layer1_node11_MUX_bit_math_h_l849_c3_c418_cond : unsigned(0 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_c418_iftrue : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_c418_iffalse : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_c418_return_output : unsigned(7 downto 0);

-- layer1_node12_MUX[bit_math_h_l860_c3_3ea5]
signal layer1_node12_MUX_bit_math_h_l860_c3_3ea5_cond : unsigned(0 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iftrue : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iffalse : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_3ea5_return_output : unsigned(7 downto 0);

-- layer1_node13_MUX[bit_math_h_l871_c3_66e4]
signal layer1_node13_MUX_bit_math_h_l871_c3_66e4_cond : unsigned(0 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_66e4_iftrue : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_66e4_iffalse : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_66e4_return_output : unsigned(7 downto 0);

-- layer1_node14_MUX[bit_math_h_l882_c3_5e4a]
signal layer1_node14_MUX_bit_math_h_l882_c3_5e4a_cond : unsigned(0 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iftrue : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iffalse : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_5e4a_return_output : unsigned(7 downto 0);

-- layer1_node15_MUX[bit_math_h_l893_c3_faee]
signal layer1_node15_MUX_bit_math_h_l893_c3_faee_cond : unsigned(0 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_faee_iftrue : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_faee_iffalse : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_faee_return_output : unsigned(7 downto 0);

-- layer1_node16_MUX[bit_math_h_l904_c3_1e1f]
signal layer1_node16_MUX_bit_math_h_l904_c3_1e1f_cond : unsigned(0 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iftrue : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iffalse : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_1e1f_return_output : unsigned(7 downto 0);

-- layer1_node17_MUX[bit_math_h_l915_c3_bbc7]
signal layer1_node17_MUX_bit_math_h_l915_c3_bbc7_cond : unsigned(0 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iftrue : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iffalse : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_bbc7_return_output : unsigned(7 downto 0);

-- layer1_node18_MUX[bit_math_h_l926_c3_15bb]
signal layer1_node18_MUX_bit_math_h_l926_c3_15bb_cond : unsigned(0 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_15bb_iftrue : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_15bb_iffalse : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_15bb_return_output : unsigned(7 downto 0);

-- layer1_node19_MUX[bit_math_h_l937_c3_3ad6]
signal layer1_node19_MUX_bit_math_h_l937_c3_3ad6_cond : unsigned(0 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iftrue : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iffalse : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_3ad6_return_output : unsigned(7 downto 0);

-- layer1_node20_MUX[bit_math_h_l948_c3_d497]
signal layer1_node20_MUX_bit_math_h_l948_c3_d497_cond : unsigned(0 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_d497_iftrue : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_d497_iffalse : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_d497_return_output : unsigned(7 downto 0);

-- layer1_node21_MUX[bit_math_h_l959_c3_0003]
signal layer1_node21_MUX_bit_math_h_l959_c3_0003_cond : unsigned(0 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_0003_iftrue : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_0003_iffalse : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_0003_return_output : unsigned(7 downto 0);

-- layer1_node22_MUX[bit_math_h_l970_c3_fb2c]
signal layer1_node22_MUX_bit_math_h_l970_c3_fb2c_cond : unsigned(0 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iftrue : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iffalse : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_fb2c_return_output : unsigned(7 downto 0);

-- layer1_node23_MUX[bit_math_h_l981_c3_c1f3]
signal layer1_node23_MUX_bit_math_h_l981_c3_c1f3_cond : unsigned(0 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iftrue : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iffalse : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_c1f3_return_output : unsigned(7 downto 0);

-- layer1_node24_MUX[bit_math_h_l992_c3_1884]
signal layer1_node24_MUX_bit_math_h_l992_c3_1884_cond : unsigned(0 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_1884_iftrue : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_1884_iffalse : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_1884_return_output : unsigned(7 downto 0);

-- layer1_node25_MUX[bit_math_h_l1003_c3_371a]
signal layer1_node25_MUX_bit_math_h_l1003_c3_371a_cond : unsigned(0 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_371a_iftrue : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_371a_iffalse : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_371a_return_output : unsigned(7 downto 0);

-- layer1_node26_MUX[bit_math_h_l1014_c3_b858]
signal layer1_node26_MUX_bit_math_h_l1014_c3_b858_cond : unsigned(0 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_b858_iftrue : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_b858_iffalse : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_b858_return_output : unsigned(7 downto 0);

-- layer1_node27_MUX[bit_math_h_l1025_c3_d07c]
signal layer1_node27_MUX_bit_math_h_l1025_c3_d07c_cond : unsigned(0 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iftrue : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iffalse : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_d07c_return_output : unsigned(7 downto 0);

-- layer1_node28_MUX[bit_math_h_l1036_c3_d560]
signal layer1_node28_MUX_bit_math_h_l1036_c3_d560_cond : unsigned(0 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_d560_iftrue : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_d560_iffalse : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_d560_return_output : unsigned(7 downto 0);

-- layer1_node29_MUX[bit_math_h_l1047_c3_9f00]
signal layer1_node29_MUX_bit_math_h_l1047_c3_9f00_cond : unsigned(0 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iftrue : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iffalse : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_9f00_return_output : unsigned(7 downto 0);

-- layer1_node30_MUX[bit_math_h_l1058_c3_e6cc]
signal layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_cond : unsigned(0 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iftrue : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iffalse : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_return_output : unsigned(7 downto 0);

-- layer1_node31_MUX[bit_math_h_l1069_c3_b1c7]
signal layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_cond : unsigned(0 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iftrue : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iffalse : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_return_output : unsigned(7 downto 0);

-- layer2_node0_MUX[bit_math_h_l1086_c3_f3d3]
signal layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iftrue : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iffalse : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_return_output : unsigned(7 downto 0);

-- layer2_node1_MUX[bit_math_h_l1097_c3_7335]
signal layer2_node1_MUX_bit_math_h_l1097_c3_7335_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_7335_iftrue : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_7335_iffalse : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_7335_return_output : unsigned(7 downto 0);

-- layer2_node2_MUX[bit_math_h_l1108_c3_bb5a]
signal layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_cond : unsigned(0 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iftrue : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iffalse : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_return_output : unsigned(7 downto 0);

-- layer2_node3_MUX[bit_math_h_l1119_c3_95be]
signal layer2_node3_MUX_bit_math_h_l1119_c3_95be_cond : unsigned(0 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_95be_iftrue : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_95be_iffalse : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_95be_return_output : unsigned(7 downto 0);

-- layer2_node4_MUX[bit_math_h_l1130_c3_0608]
signal layer2_node4_MUX_bit_math_h_l1130_c3_0608_cond : unsigned(0 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_0608_iftrue : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_0608_iffalse : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_0608_return_output : unsigned(7 downto 0);

-- layer2_node5_MUX[bit_math_h_l1141_c3_a965]
signal layer2_node5_MUX_bit_math_h_l1141_c3_a965_cond : unsigned(0 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a965_iftrue : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a965_iffalse : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_a965_return_output : unsigned(7 downto 0);

-- layer2_node6_MUX[bit_math_h_l1152_c3_be4a]
signal layer2_node6_MUX_bit_math_h_l1152_c3_be4a_cond : unsigned(0 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iftrue : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iffalse : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_be4a_return_output : unsigned(7 downto 0);

-- layer2_node7_MUX[bit_math_h_l1163_c3_4bab]
signal layer2_node7_MUX_bit_math_h_l1163_c3_4bab_cond : unsigned(0 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iftrue : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iffalse : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_4bab_return_output : unsigned(7 downto 0);

-- layer2_node8_MUX[bit_math_h_l1174_c3_24ff]
signal layer2_node8_MUX_bit_math_h_l1174_c3_24ff_cond : unsigned(0 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iftrue : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iffalse : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_24ff_return_output : unsigned(7 downto 0);

-- layer2_node9_MUX[bit_math_h_l1185_c3_e581]
signal layer2_node9_MUX_bit_math_h_l1185_c3_e581_cond : unsigned(0 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_e581_iftrue : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_e581_iffalse : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_e581_return_output : unsigned(7 downto 0);

-- layer2_node10_MUX[bit_math_h_l1196_c3_c187]
signal layer2_node10_MUX_bit_math_h_l1196_c3_c187_cond : unsigned(0 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_c187_iftrue : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_c187_iffalse : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_c187_return_output : unsigned(7 downto 0);

-- layer2_node11_MUX[bit_math_h_l1207_c3_bafc]
signal layer2_node11_MUX_bit_math_h_l1207_c3_bafc_cond : unsigned(0 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iftrue : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iffalse : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_bafc_return_output : unsigned(7 downto 0);

-- layer2_node12_MUX[bit_math_h_l1218_c3_c26f]
signal layer2_node12_MUX_bit_math_h_l1218_c3_c26f_cond : unsigned(0 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iftrue : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iffalse : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_c26f_return_output : unsigned(7 downto 0);

-- layer2_node13_MUX[bit_math_h_l1229_c3_bcb9]
signal layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_cond : unsigned(0 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iftrue : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iffalse : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_return_output : unsigned(7 downto 0);

-- layer2_node14_MUX[bit_math_h_l1240_c3_7be3]
signal layer2_node14_MUX_bit_math_h_l1240_c3_7be3_cond : unsigned(0 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iftrue : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iffalse : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_7be3_return_output : unsigned(7 downto 0);

-- layer2_node15_MUX[bit_math_h_l1251_c3_1e63]
signal layer2_node15_MUX_bit_math_h_l1251_c3_1e63_cond : unsigned(0 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iftrue : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iffalse : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_1e63_return_output : unsigned(7 downto 0);

-- layer3_node0_MUX[bit_math_h_l1268_c3_e356]
signal layer3_node0_MUX_bit_math_h_l1268_c3_e356_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_e356_iftrue : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_e356_iffalse : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_e356_return_output : unsigned(7 downto 0);

-- layer3_node1_MUX[bit_math_h_l1279_c3_3873]
signal layer3_node1_MUX_bit_math_h_l1279_c3_3873_cond : unsigned(0 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_3873_iftrue : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_3873_iffalse : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_3873_return_output : unsigned(7 downto 0);

-- layer3_node2_MUX[bit_math_h_l1290_c3_4ec7]
signal layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_cond : unsigned(0 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iftrue : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iffalse : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_return_output : unsigned(7 downto 0);

-- layer3_node3_MUX[bit_math_h_l1301_c3_29f9]
signal layer3_node3_MUX_bit_math_h_l1301_c3_29f9_cond : unsigned(0 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iftrue : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iffalse : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_29f9_return_output : unsigned(7 downto 0);

-- layer3_node4_MUX[bit_math_h_l1312_c3_b484]
signal layer3_node4_MUX_bit_math_h_l1312_c3_b484_cond : unsigned(0 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_b484_iftrue : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_b484_iffalse : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_b484_return_output : unsigned(7 downto 0);

-- layer3_node5_MUX[bit_math_h_l1323_c3_e63b]
signal layer3_node5_MUX_bit_math_h_l1323_c3_e63b_cond : unsigned(0 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iftrue : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iffalse : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_e63b_return_output : unsigned(7 downto 0);

-- layer3_node6_MUX[bit_math_h_l1334_c3_5def]
signal layer3_node6_MUX_bit_math_h_l1334_c3_5def_cond : unsigned(0 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_5def_iftrue : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_5def_iffalse : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_5def_return_output : unsigned(7 downto 0);

-- layer3_node7_MUX[bit_math_h_l1345_c3_3cb2]
signal layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_cond : unsigned(0 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iftrue : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iffalse : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_return_output : unsigned(7 downto 0);

-- layer4_node0_MUX[bit_math_h_l1362_c3_fa41]
signal layer4_node0_MUX_bit_math_h_l1362_c3_fa41_cond : unsigned(0 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iftrue : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iffalse : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_fa41_return_output : unsigned(7 downto 0);

-- layer4_node1_MUX[bit_math_h_l1373_c3_223f]
signal layer4_node1_MUX_bit_math_h_l1373_c3_223f_cond : unsigned(0 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_223f_iftrue : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_223f_iffalse : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_223f_return_output : unsigned(7 downto 0);

-- layer4_node2_MUX[bit_math_h_l1384_c3_470b]
signal layer4_node2_MUX_bit_math_h_l1384_c3_470b_cond : unsigned(0 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_470b_iftrue : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_470b_iffalse : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_470b_return_output : unsigned(7 downto 0);

-- layer4_node3_MUX[bit_math_h_l1395_c3_68f4]
signal layer4_node3_MUX_bit_math_h_l1395_c3_68f4_cond : unsigned(0 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iftrue : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iffalse : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_68f4_return_output : unsigned(7 downto 0);

-- layer5_node0_MUX[bit_math_h_l1412_c3_e3bb]
signal layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_cond : unsigned(0 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iftrue : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iffalse : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_return_output : unsigned(7 downto 0);

-- layer5_node1_MUX[bit_math_h_l1423_c3_47e8]
signal layer5_node1_MUX_bit_math_h_l1423_c3_47e8_cond : unsigned(0 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iftrue : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iffalse : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_47e8_return_output : unsigned(7 downto 0);

-- layer6_node0_MUX[bit_math_h_l1440_c3_7682]
signal layer6_node0_MUX_bit_math_h_l1440_c3_7682_cond : unsigned(0 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_7682_iftrue : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_7682_iffalse : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_7682_return_output : unsigned(7 downto 0);

function uint7_0_0( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint7_1_1( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint7_2_2( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint7_3_3( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;

function uint7_4_4( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(4- i);
      end loop;
return return_output;
end function;

function uint7_5_5( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(5- i);
      end loop;
return return_output;
end function;

function uint7_6_6( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(6- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_70c7
layer0_node0_MUX_bit_math_h_l18_c3_70c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_70c7_cond,
layer0_node0_MUX_bit_math_h_l18_c3_70c7_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_70c7_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_70c7_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_dc12
layer0_node1_MUX_bit_math_h_l29_c3_dc12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_dc12_cond,
layer0_node1_MUX_bit_math_h_l29_c3_dc12_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_dc12_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_dc12_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_3404
layer0_node2_MUX_bit_math_h_l40_c3_3404 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_3404_cond,
layer0_node2_MUX_bit_math_h_l40_c3_3404_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_3404_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_3404_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_cc01
layer0_node3_MUX_bit_math_h_l51_c3_cc01 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_cc01_cond,
layer0_node3_MUX_bit_math_h_l51_c3_cc01_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_cc01_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_cc01_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_7793
layer0_node4_MUX_bit_math_h_l62_c3_7793 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_7793_cond,
layer0_node4_MUX_bit_math_h_l62_c3_7793_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_7793_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_7793_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_2acd
layer0_node5_MUX_bit_math_h_l73_c3_2acd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_2acd_cond,
layer0_node5_MUX_bit_math_h_l73_c3_2acd_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_2acd_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_2acd_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_494b
layer0_node6_MUX_bit_math_h_l84_c3_494b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_494b_cond,
layer0_node6_MUX_bit_math_h_l84_c3_494b_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_494b_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_494b_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_daab
layer0_node7_MUX_bit_math_h_l95_c3_daab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_daab_cond,
layer0_node7_MUX_bit_math_h_l95_c3_daab_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_daab_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_daab_return_output);

-- layer0_node8_MUX_bit_math_h_l106_c3_d50d
layer0_node8_MUX_bit_math_h_l106_c3_d50d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node8_MUX_bit_math_h_l106_c3_d50d_cond,
layer0_node8_MUX_bit_math_h_l106_c3_d50d_iftrue,
layer0_node8_MUX_bit_math_h_l106_c3_d50d_iffalse,
layer0_node8_MUX_bit_math_h_l106_c3_d50d_return_output);

-- layer0_node9_MUX_bit_math_h_l117_c3_c9ee
layer0_node9_MUX_bit_math_h_l117_c3_c9ee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node9_MUX_bit_math_h_l117_c3_c9ee_cond,
layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iftrue,
layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iffalse,
layer0_node9_MUX_bit_math_h_l117_c3_c9ee_return_output);

-- layer0_node10_MUX_bit_math_h_l128_c3_06d1
layer0_node10_MUX_bit_math_h_l128_c3_06d1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node10_MUX_bit_math_h_l128_c3_06d1_cond,
layer0_node10_MUX_bit_math_h_l128_c3_06d1_iftrue,
layer0_node10_MUX_bit_math_h_l128_c3_06d1_iffalse,
layer0_node10_MUX_bit_math_h_l128_c3_06d1_return_output);

-- layer0_node11_MUX_bit_math_h_l139_c3_13dc
layer0_node11_MUX_bit_math_h_l139_c3_13dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node11_MUX_bit_math_h_l139_c3_13dc_cond,
layer0_node11_MUX_bit_math_h_l139_c3_13dc_iftrue,
layer0_node11_MUX_bit_math_h_l139_c3_13dc_iffalse,
layer0_node11_MUX_bit_math_h_l139_c3_13dc_return_output);

-- layer0_node12_MUX_bit_math_h_l150_c3_af2c
layer0_node12_MUX_bit_math_h_l150_c3_af2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node12_MUX_bit_math_h_l150_c3_af2c_cond,
layer0_node12_MUX_bit_math_h_l150_c3_af2c_iftrue,
layer0_node12_MUX_bit_math_h_l150_c3_af2c_iffalse,
layer0_node12_MUX_bit_math_h_l150_c3_af2c_return_output);

-- layer0_node13_MUX_bit_math_h_l161_c3_c865
layer0_node13_MUX_bit_math_h_l161_c3_c865 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node13_MUX_bit_math_h_l161_c3_c865_cond,
layer0_node13_MUX_bit_math_h_l161_c3_c865_iftrue,
layer0_node13_MUX_bit_math_h_l161_c3_c865_iffalse,
layer0_node13_MUX_bit_math_h_l161_c3_c865_return_output);

-- layer0_node14_MUX_bit_math_h_l172_c3_1937
layer0_node14_MUX_bit_math_h_l172_c3_1937 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node14_MUX_bit_math_h_l172_c3_1937_cond,
layer0_node14_MUX_bit_math_h_l172_c3_1937_iftrue,
layer0_node14_MUX_bit_math_h_l172_c3_1937_iffalse,
layer0_node14_MUX_bit_math_h_l172_c3_1937_return_output);

-- layer0_node15_MUX_bit_math_h_l183_c3_6211
layer0_node15_MUX_bit_math_h_l183_c3_6211 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node15_MUX_bit_math_h_l183_c3_6211_cond,
layer0_node15_MUX_bit_math_h_l183_c3_6211_iftrue,
layer0_node15_MUX_bit_math_h_l183_c3_6211_iffalse,
layer0_node15_MUX_bit_math_h_l183_c3_6211_return_output);

-- layer0_node16_MUX_bit_math_h_l194_c3_6e24
layer0_node16_MUX_bit_math_h_l194_c3_6e24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node16_MUX_bit_math_h_l194_c3_6e24_cond,
layer0_node16_MUX_bit_math_h_l194_c3_6e24_iftrue,
layer0_node16_MUX_bit_math_h_l194_c3_6e24_iffalse,
layer0_node16_MUX_bit_math_h_l194_c3_6e24_return_output);

-- layer0_node17_MUX_bit_math_h_l205_c3_4b2c
layer0_node17_MUX_bit_math_h_l205_c3_4b2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node17_MUX_bit_math_h_l205_c3_4b2c_cond,
layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iftrue,
layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iffalse,
layer0_node17_MUX_bit_math_h_l205_c3_4b2c_return_output);

-- layer0_node18_MUX_bit_math_h_l216_c3_0b83
layer0_node18_MUX_bit_math_h_l216_c3_0b83 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node18_MUX_bit_math_h_l216_c3_0b83_cond,
layer0_node18_MUX_bit_math_h_l216_c3_0b83_iftrue,
layer0_node18_MUX_bit_math_h_l216_c3_0b83_iffalse,
layer0_node18_MUX_bit_math_h_l216_c3_0b83_return_output);

-- layer0_node19_MUX_bit_math_h_l227_c3_1e36
layer0_node19_MUX_bit_math_h_l227_c3_1e36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node19_MUX_bit_math_h_l227_c3_1e36_cond,
layer0_node19_MUX_bit_math_h_l227_c3_1e36_iftrue,
layer0_node19_MUX_bit_math_h_l227_c3_1e36_iffalse,
layer0_node19_MUX_bit_math_h_l227_c3_1e36_return_output);

-- layer0_node20_MUX_bit_math_h_l238_c3_5458
layer0_node20_MUX_bit_math_h_l238_c3_5458 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node20_MUX_bit_math_h_l238_c3_5458_cond,
layer0_node20_MUX_bit_math_h_l238_c3_5458_iftrue,
layer0_node20_MUX_bit_math_h_l238_c3_5458_iffalse,
layer0_node20_MUX_bit_math_h_l238_c3_5458_return_output);

-- layer0_node21_MUX_bit_math_h_l249_c3_c173
layer0_node21_MUX_bit_math_h_l249_c3_c173 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node21_MUX_bit_math_h_l249_c3_c173_cond,
layer0_node21_MUX_bit_math_h_l249_c3_c173_iftrue,
layer0_node21_MUX_bit_math_h_l249_c3_c173_iffalse,
layer0_node21_MUX_bit_math_h_l249_c3_c173_return_output);

-- layer0_node22_MUX_bit_math_h_l260_c3_fce5
layer0_node22_MUX_bit_math_h_l260_c3_fce5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node22_MUX_bit_math_h_l260_c3_fce5_cond,
layer0_node22_MUX_bit_math_h_l260_c3_fce5_iftrue,
layer0_node22_MUX_bit_math_h_l260_c3_fce5_iffalse,
layer0_node22_MUX_bit_math_h_l260_c3_fce5_return_output);

-- layer0_node23_MUX_bit_math_h_l271_c3_a82d
layer0_node23_MUX_bit_math_h_l271_c3_a82d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node23_MUX_bit_math_h_l271_c3_a82d_cond,
layer0_node23_MUX_bit_math_h_l271_c3_a82d_iftrue,
layer0_node23_MUX_bit_math_h_l271_c3_a82d_iffalse,
layer0_node23_MUX_bit_math_h_l271_c3_a82d_return_output);

-- layer0_node24_MUX_bit_math_h_l282_c3_6611
layer0_node24_MUX_bit_math_h_l282_c3_6611 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node24_MUX_bit_math_h_l282_c3_6611_cond,
layer0_node24_MUX_bit_math_h_l282_c3_6611_iftrue,
layer0_node24_MUX_bit_math_h_l282_c3_6611_iffalse,
layer0_node24_MUX_bit_math_h_l282_c3_6611_return_output);

-- layer0_node25_MUX_bit_math_h_l293_c3_b4b9
layer0_node25_MUX_bit_math_h_l293_c3_b4b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node25_MUX_bit_math_h_l293_c3_b4b9_cond,
layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iftrue,
layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iffalse,
layer0_node25_MUX_bit_math_h_l293_c3_b4b9_return_output);

-- layer0_node26_MUX_bit_math_h_l304_c3_2bce
layer0_node26_MUX_bit_math_h_l304_c3_2bce : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node26_MUX_bit_math_h_l304_c3_2bce_cond,
layer0_node26_MUX_bit_math_h_l304_c3_2bce_iftrue,
layer0_node26_MUX_bit_math_h_l304_c3_2bce_iffalse,
layer0_node26_MUX_bit_math_h_l304_c3_2bce_return_output);

-- layer0_node27_MUX_bit_math_h_l315_c3_7789
layer0_node27_MUX_bit_math_h_l315_c3_7789 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node27_MUX_bit_math_h_l315_c3_7789_cond,
layer0_node27_MUX_bit_math_h_l315_c3_7789_iftrue,
layer0_node27_MUX_bit_math_h_l315_c3_7789_iffalse,
layer0_node27_MUX_bit_math_h_l315_c3_7789_return_output);

-- layer0_node28_MUX_bit_math_h_l326_c3_098d
layer0_node28_MUX_bit_math_h_l326_c3_098d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node28_MUX_bit_math_h_l326_c3_098d_cond,
layer0_node28_MUX_bit_math_h_l326_c3_098d_iftrue,
layer0_node28_MUX_bit_math_h_l326_c3_098d_iffalse,
layer0_node28_MUX_bit_math_h_l326_c3_098d_return_output);

-- layer0_node29_MUX_bit_math_h_l337_c3_9c87
layer0_node29_MUX_bit_math_h_l337_c3_9c87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node29_MUX_bit_math_h_l337_c3_9c87_cond,
layer0_node29_MUX_bit_math_h_l337_c3_9c87_iftrue,
layer0_node29_MUX_bit_math_h_l337_c3_9c87_iffalse,
layer0_node29_MUX_bit_math_h_l337_c3_9c87_return_output);

-- layer0_node30_MUX_bit_math_h_l348_c3_6b0d
layer0_node30_MUX_bit_math_h_l348_c3_6b0d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node30_MUX_bit_math_h_l348_c3_6b0d_cond,
layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iftrue,
layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iffalse,
layer0_node30_MUX_bit_math_h_l348_c3_6b0d_return_output);

-- layer0_node31_MUX_bit_math_h_l359_c3_5065
layer0_node31_MUX_bit_math_h_l359_c3_5065 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node31_MUX_bit_math_h_l359_c3_5065_cond,
layer0_node31_MUX_bit_math_h_l359_c3_5065_iftrue,
layer0_node31_MUX_bit_math_h_l359_c3_5065_iffalse,
layer0_node31_MUX_bit_math_h_l359_c3_5065_return_output);

-- layer0_node32_MUX_bit_math_h_l370_c3_4893
layer0_node32_MUX_bit_math_h_l370_c3_4893 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node32_MUX_bit_math_h_l370_c3_4893_cond,
layer0_node32_MUX_bit_math_h_l370_c3_4893_iftrue,
layer0_node32_MUX_bit_math_h_l370_c3_4893_iffalse,
layer0_node32_MUX_bit_math_h_l370_c3_4893_return_output);

-- layer0_node33_MUX_bit_math_h_l381_c3_8132
layer0_node33_MUX_bit_math_h_l381_c3_8132 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node33_MUX_bit_math_h_l381_c3_8132_cond,
layer0_node33_MUX_bit_math_h_l381_c3_8132_iftrue,
layer0_node33_MUX_bit_math_h_l381_c3_8132_iffalse,
layer0_node33_MUX_bit_math_h_l381_c3_8132_return_output);

-- layer0_node34_MUX_bit_math_h_l392_c3_59bd
layer0_node34_MUX_bit_math_h_l392_c3_59bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node34_MUX_bit_math_h_l392_c3_59bd_cond,
layer0_node34_MUX_bit_math_h_l392_c3_59bd_iftrue,
layer0_node34_MUX_bit_math_h_l392_c3_59bd_iffalse,
layer0_node34_MUX_bit_math_h_l392_c3_59bd_return_output);

-- layer0_node35_MUX_bit_math_h_l403_c3_6326
layer0_node35_MUX_bit_math_h_l403_c3_6326 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node35_MUX_bit_math_h_l403_c3_6326_cond,
layer0_node35_MUX_bit_math_h_l403_c3_6326_iftrue,
layer0_node35_MUX_bit_math_h_l403_c3_6326_iffalse,
layer0_node35_MUX_bit_math_h_l403_c3_6326_return_output);

-- layer0_node36_MUX_bit_math_h_l414_c3_7348
layer0_node36_MUX_bit_math_h_l414_c3_7348 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node36_MUX_bit_math_h_l414_c3_7348_cond,
layer0_node36_MUX_bit_math_h_l414_c3_7348_iftrue,
layer0_node36_MUX_bit_math_h_l414_c3_7348_iffalse,
layer0_node36_MUX_bit_math_h_l414_c3_7348_return_output);

-- layer0_node37_MUX_bit_math_h_l425_c3_f929
layer0_node37_MUX_bit_math_h_l425_c3_f929 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node37_MUX_bit_math_h_l425_c3_f929_cond,
layer0_node37_MUX_bit_math_h_l425_c3_f929_iftrue,
layer0_node37_MUX_bit_math_h_l425_c3_f929_iffalse,
layer0_node37_MUX_bit_math_h_l425_c3_f929_return_output);

-- layer0_node38_MUX_bit_math_h_l436_c3_d3a0
layer0_node38_MUX_bit_math_h_l436_c3_d3a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node38_MUX_bit_math_h_l436_c3_d3a0_cond,
layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iftrue,
layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iffalse,
layer0_node38_MUX_bit_math_h_l436_c3_d3a0_return_output);

-- layer0_node39_MUX_bit_math_h_l447_c3_7b35
layer0_node39_MUX_bit_math_h_l447_c3_7b35 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node39_MUX_bit_math_h_l447_c3_7b35_cond,
layer0_node39_MUX_bit_math_h_l447_c3_7b35_iftrue,
layer0_node39_MUX_bit_math_h_l447_c3_7b35_iffalse,
layer0_node39_MUX_bit_math_h_l447_c3_7b35_return_output);

-- layer0_node40_MUX_bit_math_h_l458_c3_426b
layer0_node40_MUX_bit_math_h_l458_c3_426b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node40_MUX_bit_math_h_l458_c3_426b_cond,
layer0_node40_MUX_bit_math_h_l458_c3_426b_iftrue,
layer0_node40_MUX_bit_math_h_l458_c3_426b_iffalse,
layer0_node40_MUX_bit_math_h_l458_c3_426b_return_output);

-- layer0_node41_MUX_bit_math_h_l469_c3_47d5
layer0_node41_MUX_bit_math_h_l469_c3_47d5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node41_MUX_bit_math_h_l469_c3_47d5_cond,
layer0_node41_MUX_bit_math_h_l469_c3_47d5_iftrue,
layer0_node41_MUX_bit_math_h_l469_c3_47d5_iffalse,
layer0_node41_MUX_bit_math_h_l469_c3_47d5_return_output);

-- layer0_node42_MUX_bit_math_h_l480_c3_50c3
layer0_node42_MUX_bit_math_h_l480_c3_50c3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node42_MUX_bit_math_h_l480_c3_50c3_cond,
layer0_node42_MUX_bit_math_h_l480_c3_50c3_iftrue,
layer0_node42_MUX_bit_math_h_l480_c3_50c3_iffalse,
layer0_node42_MUX_bit_math_h_l480_c3_50c3_return_output);

-- layer0_node43_MUX_bit_math_h_l491_c3_6ed7
layer0_node43_MUX_bit_math_h_l491_c3_6ed7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node43_MUX_bit_math_h_l491_c3_6ed7_cond,
layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iftrue,
layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iffalse,
layer0_node43_MUX_bit_math_h_l491_c3_6ed7_return_output);

-- layer0_node44_MUX_bit_math_h_l502_c3_84a4
layer0_node44_MUX_bit_math_h_l502_c3_84a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node44_MUX_bit_math_h_l502_c3_84a4_cond,
layer0_node44_MUX_bit_math_h_l502_c3_84a4_iftrue,
layer0_node44_MUX_bit_math_h_l502_c3_84a4_iffalse,
layer0_node44_MUX_bit_math_h_l502_c3_84a4_return_output);

-- layer0_node45_MUX_bit_math_h_l513_c3_552e
layer0_node45_MUX_bit_math_h_l513_c3_552e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node45_MUX_bit_math_h_l513_c3_552e_cond,
layer0_node45_MUX_bit_math_h_l513_c3_552e_iftrue,
layer0_node45_MUX_bit_math_h_l513_c3_552e_iffalse,
layer0_node45_MUX_bit_math_h_l513_c3_552e_return_output);

-- layer0_node46_MUX_bit_math_h_l524_c3_42cd
layer0_node46_MUX_bit_math_h_l524_c3_42cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node46_MUX_bit_math_h_l524_c3_42cd_cond,
layer0_node46_MUX_bit_math_h_l524_c3_42cd_iftrue,
layer0_node46_MUX_bit_math_h_l524_c3_42cd_iffalse,
layer0_node46_MUX_bit_math_h_l524_c3_42cd_return_output);

-- layer0_node47_MUX_bit_math_h_l535_c3_18b2
layer0_node47_MUX_bit_math_h_l535_c3_18b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node47_MUX_bit_math_h_l535_c3_18b2_cond,
layer0_node47_MUX_bit_math_h_l535_c3_18b2_iftrue,
layer0_node47_MUX_bit_math_h_l535_c3_18b2_iffalse,
layer0_node47_MUX_bit_math_h_l535_c3_18b2_return_output);

-- layer0_node48_MUX_bit_math_h_l546_c3_e9fe
layer0_node48_MUX_bit_math_h_l546_c3_e9fe : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node48_MUX_bit_math_h_l546_c3_e9fe_cond,
layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iftrue,
layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iffalse,
layer0_node48_MUX_bit_math_h_l546_c3_e9fe_return_output);

-- layer0_node49_MUX_bit_math_h_l557_c3_68c1
layer0_node49_MUX_bit_math_h_l557_c3_68c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node49_MUX_bit_math_h_l557_c3_68c1_cond,
layer0_node49_MUX_bit_math_h_l557_c3_68c1_iftrue,
layer0_node49_MUX_bit_math_h_l557_c3_68c1_iffalse,
layer0_node49_MUX_bit_math_h_l557_c3_68c1_return_output);

-- layer0_node50_MUX_bit_math_h_l568_c3_8ec7
layer0_node50_MUX_bit_math_h_l568_c3_8ec7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node50_MUX_bit_math_h_l568_c3_8ec7_cond,
layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iftrue,
layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iffalse,
layer0_node50_MUX_bit_math_h_l568_c3_8ec7_return_output);

-- layer0_node51_MUX_bit_math_h_l579_c3_5985
layer0_node51_MUX_bit_math_h_l579_c3_5985 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node51_MUX_bit_math_h_l579_c3_5985_cond,
layer0_node51_MUX_bit_math_h_l579_c3_5985_iftrue,
layer0_node51_MUX_bit_math_h_l579_c3_5985_iffalse,
layer0_node51_MUX_bit_math_h_l579_c3_5985_return_output);

-- layer0_node52_MUX_bit_math_h_l590_c3_90c2
layer0_node52_MUX_bit_math_h_l590_c3_90c2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node52_MUX_bit_math_h_l590_c3_90c2_cond,
layer0_node52_MUX_bit_math_h_l590_c3_90c2_iftrue,
layer0_node52_MUX_bit_math_h_l590_c3_90c2_iffalse,
layer0_node52_MUX_bit_math_h_l590_c3_90c2_return_output);

-- layer0_node53_MUX_bit_math_h_l601_c3_5a9e
layer0_node53_MUX_bit_math_h_l601_c3_5a9e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node53_MUX_bit_math_h_l601_c3_5a9e_cond,
layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iftrue,
layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iffalse,
layer0_node53_MUX_bit_math_h_l601_c3_5a9e_return_output);

-- layer0_node54_MUX_bit_math_h_l612_c3_235a
layer0_node54_MUX_bit_math_h_l612_c3_235a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node54_MUX_bit_math_h_l612_c3_235a_cond,
layer0_node54_MUX_bit_math_h_l612_c3_235a_iftrue,
layer0_node54_MUX_bit_math_h_l612_c3_235a_iffalse,
layer0_node54_MUX_bit_math_h_l612_c3_235a_return_output);

-- layer0_node55_MUX_bit_math_h_l623_c3_1dea
layer0_node55_MUX_bit_math_h_l623_c3_1dea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node55_MUX_bit_math_h_l623_c3_1dea_cond,
layer0_node55_MUX_bit_math_h_l623_c3_1dea_iftrue,
layer0_node55_MUX_bit_math_h_l623_c3_1dea_iffalse,
layer0_node55_MUX_bit_math_h_l623_c3_1dea_return_output);

-- layer0_node56_MUX_bit_math_h_l634_c3_f6e3
layer0_node56_MUX_bit_math_h_l634_c3_f6e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node56_MUX_bit_math_h_l634_c3_f6e3_cond,
layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iftrue,
layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iffalse,
layer0_node56_MUX_bit_math_h_l634_c3_f6e3_return_output);

-- layer0_node57_MUX_bit_math_h_l645_c3_eeb0
layer0_node57_MUX_bit_math_h_l645_c3_eeb0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node57_MUX_bit_math_h_l645_c3_eeb0_cond,
layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iftrue,
layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iffalse,
layer0_node57_MUX_bit_math_h_l645_c3_eeb0_return_output);

-- layer0_node58_MUX_bit_math_h_l656_c3_b995
layer0_node58_MUX_bit_math_h_l656_c3_b995 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node58_MUX_bit_math_h_l656_c3_b995_cond,
layer0_node58_MUX_bit_math_h_l656_c3_b995_iftrue,
layer0_node58_MUX_bit_math_h_l656_c3_b995_iffalse,
layer0_node58_MUX_bit_math_h_l656_c3_b995_return_output);

-- layer0_node59_MUX_bit_math_h_l667_c3_b104
layer0_node59_MUX_bit_math_h_l667_c3_b104 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node59_MUX_bit_math_h_l667_c3_b104_cond,
layer0_node59_MUX_bit_math_h_l667_c3_b104_iftrue,
layer0_node59_MUX_bit_math_h_l667_c3_b104_iffalse,
layer0_node59_MUX_bit_math_h_l667_c3_b104_return_output);

-- layer0_node60_MUX_bit_math_h_l678_c3_7571
layer0_node60_MUX_bit_math_h_l678_c3_7571 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node60_MUX_bit_math_h_l678_c3_7571_cond,
layer0_node60_MUX_bit_math_h_l678_c3_7571_iftrue,
layer0_node60_MUX_bit_math_h_l678_c3_7571_iffalse,
layer0_node60_MUX_bit_math_h_l678_c3_7571_return_output);

-- layer0_node61_MUX_bit_math_h_l689_c3_580e
layer0_node61_MUX_bit_math_h_l689_c3_580e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node61_MUX_bit_math_h_l689_c3_580e_cond,
layer0_node61_MUX_bit_math_h_l689_c3_580e_iftrue,
layer0_node61_MUX_bit_math_h_l689_c3_580e_iffalse,
layer0_node61_MUX_bit_math_h_l689_c3_580e_return_output);

-- layer0_node62_MUX_bit_math_h_l700_c3_9f5f
layer0_node62_MUX_bit_math_h_l700_c3_9f5f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node62_MUX_bit_math_h_l700_c3_9f5f_cond,
layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iftrue,
layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iffalse,
layer0_node62_MUX_bit_math_h_l700_c3_9f5f_return_output);

-- layer0_node63_MUX_bit_math_h_l711_c3_17f2
layer0_node63_MUX_bit_math_h_l711_c3_17f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node63_MUX_bit_math_h_l711_c3_17f2_cond,
layer0_node63_MUX_bit_math_h_l711_c3_17f2_iftrue,
layer0_node63_MUX_bit_math_h_l711_c3_17f2_iffalse,
layer0_node63_MUX_bit_math_h_l711_c3_17f2_return_output);

-- layer1_node0_MUX_bit_math_h_l728_c3_23e3
layer1_node0_MUX_bit_math_h_l728_c3_23e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l728_c3_23e3_cond,
layer1_node0_MUX_bit_math_h_l728_c3_23e3_iftrue,
layer1_node0_MUX_bit_math_h_l728_c3_23e3_iffalse,
layer1_node0_MUX_bit_math_h_l728_c3_23e3_return_output);

-- layer1_node1_MUX_bit_math_h_l739_c3_57f6
layer1_node1_MUX_bit_math_h_l739_c3_57f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l739_c3_57f6_cond,
layer1_node1_MUX_bit_math_h_l739_c3_57f6_iftrue,
layer1_node1_MUX_bit_math_h_l739_c3_57f6_iffalse,
layer1_node1_MUX_bit_math_h_l739_c3_57f6_return_output);

-- layer1_node2_MUX_bit_math_h_l750_c3_b86b
layer1_node2_MUX_bit_math_h_l750_c3_b86b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l750_c3_b86b_cond,
layer1_node2_MUX_bit_math_h_l750_c3_b86b_iftrue,
layer1_node2_MUX_bit_math_h_l750_c3_b86b_iffalse,
layer1_node2_MUX_bit_math_h_l750_c3_b86b_return_output);

-- layer1_node3_MUX_bit_math_h_l761_c3_2586
layer1_node3_MUX_bit_math_h_l761_c3_2586 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l761_c3_2586_cond,
layer1_node3_MUX_bit_math_h_l761_c3_2586_iftrue,
layer1_node3_MUX_bit_math_h_l761_c3_2586_iffalse,
layer1_node3_MUX_bit_math_h_l761_c3_2586_return_output);

-- layer1_node4_MUX_bit_math_h_l772_c3_857f
layer1_node4_MUX_bit_math_h_l772_c3_857f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node4_MUX_bit_math_h_l772_c3_857f_cond,
layer1_node4_MUX_bit_math_h_l772_c3_857f_iftrue,
layer1_node4_MUX_bit_math_h_l772_c3_857f_iffalse,
layer1_node4_MUX_bit_math_h_l772_c3_857f_return_output);

-- layer1_node5_MUX_bit_math_h_l783_c3_f8bc
layer1_node5_MUX_bit_math_h_l783_c3_f8bc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node5_MUX_bit_math_h_l783_c3_f8bc_cond,
layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iftrue,
layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iffalse,
layer1_node5_MUX_bit_math_h_l783_c3_f8bc_return_output);

-- layer1_node6_MUX_bit_math_h_l794_c3_f4dd
layer1_node6_MUX_bit_math_h_l794_c3_f4dd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node6_MUX_bit_math_h_l794_c3_f4dd_cond,
layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iftrue,
layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iffalse,
layer1_node6_MUX_bit_math_h_l794_c3_f4dd_return_output);

-- layer1_node7_MUX_bit_math_h_l805_c3_e535
layer1_node7_MUX_bit_math_h_l805_c3_e535 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node7_MUX_bit_math_h_l805_c3_e535_cond,
layer1_node7_MUX_bit_math_h_l805_c3_e535_iftrue,
layer1_node7_MUX_bit_math_h_l805_c3_e535_iffalse,
layer1_node7_MUX_bit_math_h_l805_c3_e535_return_output);

-- layer1_node8_MUX_bit_math_h_l816_c3_e51d
layer1_node8_MUX_bit_math_h_l816_c3_e51d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node8_MUX_bit_math_h_l816_c3_e51d_cond,
layer1_node8_MUX_bit_math_h_l816_c3_e51d_iftrue,
layer1_node8_MUX_bit_math_h_l816_c3_e51d_iffalse,
layer1_node8_MUX_bit_math_h_l816_c3_e51d_return_output);

-- layer1_node9_MUX_bit_math_h_l827_c3_4f17
layer1_node9_MUX_bit_math_h_l827_c3_4f17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node9_MUX_bit_math_h_l827_c3_4f17_cond,
layer1_node9_MUX_bit_math_h_l827_c3_4f17_iftrue,
layer1_node9_MUX_bit_math_h_l827_c3_4f17_iffalse,
layer1_node9_MUX_bit_math_h_l827_c3_4f17_return_output);

-- layer1_node10_MUX_bit_math_h_l838_c3_8caa
layer1_node10_MUX_bit_math_h_l838_c3_8caa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node10_MUX_bit_math_h_l838_c3_8caa_cond,
layer1_node10_MUX_bit_math_h_l838_c3_8caa_iftrue,
layer1_node10_MUX_bit_math_h_l838_c3_8caa_iffalse,
layer1_node10_MUX_bit_math_h_l838_c3_8caa_return_output);

-- layer1_node11_MUX_bit_math_h_l849_c3_c418
layer1_node11_MUX_bit_math_h_l849_c3_c418 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node11_MUX_bit_math_h_l849_c3_c418_cond,
layer1_node11_MUX_bit_math_h_l849_c3_c418_iftrue,
layer1_node11_MUX_bit_math_h_l849_c3_c418_iffalse,
layer1_node11_MUX_bit_math_h_l849_c3_c418_return_output);

-- layer1_node12_MUX_bit_math_h_l860_c3_3ea5
layer1_node12_MUX_bit_math_h_l860_c3_3ea5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node12_MUX_bit_math_h_l860_c3_3ea5_cond,
layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iftrue,
layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iffalse,
layer1_node12_MUX_bit_math_h_l860_c3_3ea5_return_output);

-- layer1_node13_MUX_bit_math_h_l871_c3_66e4
layer1_node13_MUX_bit_math_h_l871_c3_66e4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node13_MUX_bit_math_h_l871_c3_66e4_cond,
layer1_node13_MUX_bit_math_h_l871_c3_66e4_iftrue,
layer1_node13_MUX_bit_math_h_l871_c3_66e4_iffalse,
layer1_node13_MUX_bit_math_h_l871_c3_66e4_return_output);

-- layer1_node14_MUX_bit_math_h_l882_c3_5e4a
layer1_node14_MUX_bit_math_h_l882_c3_5e4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node14_MUX_bit_math_h_l882_c3_5e4a_cond,
layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iftrue,
layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iffalse,
layer1_node14_MUX_bit_math_h_l882_c3_5e4a_return_output);

-- layer1_node15_MUX_bit_math_h_l893_c3_faee
layer1_node15_MUX_bit_math_h_l893_c3_faee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node15_MUX_bit_math_h_l893_c3_faee_cond,
layer1_node15_MUX_bit_math_h_l893_c3_faee_iftrue,
layer1_node15_MUX_bit_math_h_l893_c3_faee_iffalse,
layer1_node15_MUX_bit_math_h_l893_c3_faee_return_output);

-- layer1_node16_MUX_bit_math_h_l904_c3_1e1f
layer1_node16_MUX_bit_math_h_l904_c3_1e1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node16_MUX_bit_math_h_l904_c3_1e1f_cond,
layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iftrue,
layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iffalse,
layer1_node16_MUX_bit_math_h_l904_c3_1e1f_return_output);

-- layer1_node17_MUX_bit_math_h_l915_c3_bbc7
layer1_node17_MUX_bit_math_h_l915_c3_bbc7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node17_MUX_bit_math_h_l915_c3_bbc7_cond,
layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iftrue,
layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iffalse,
layer1_node17_MUX_bit_math_h_l915_c3_bbc7_return_output);

-- layer1_node18_MUX_bit_math_h_l926_c3_15bb
layer1_node18_MUX_bit_math_h_l926_c3_15bb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node18_MUX_bit_math_h_l926_c3_15bb_cond,
layer1_node18_MUX_bit_math_h_l926_c3_15bb_iftrue,
layer1_node18_MUX_bit_math_h_l926_c3_15bb_iffalse,
layer1_node18_MUX_bit_math_h_l926_c3_15bb_return_output);

-- layer1_node19_MUX_bit_math_h_l937_c3_3ad6
layer1_node19_MUX_bit_math_h_l937_c3_3ad6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node19_MUX_bit_math_h_l937_c3_3ad6_cond,
layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iftrue,
layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iffalse,
layer1_node19_MUX_bit_math_h_l937_c3_3ad6_return_output);

-- layer1_node20_MUX_bit_math_h_l948_c3_d497
layer1_node20_MUX_bit_math_h_l948_c3_d497 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node20_MUX_bit_math_h_l948_c3_d497_cond,
layer1_node20_MUX_bit_math_h_l948_c3_d497_iftrue,
layer1_node20_MUX_bit_math_h_l948_c3_d497_iffalse,
layer1_node20_MUX_bit_math_h_l948_c3_d497_return_output);

-- layer1_node21_MUX_bit_math_h_l959_c3_0003
layer1_node21_MUX_bit_math_h_l959_c3_0003 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node21_MUX_bit_math_h_l959_c3_0003_cond,
layer1_node21_MUX_bit_math_h_l959_c3_0003_iftrue,
layer1_node21_MUX_bit_math_h_l959_c3_0003_iffalse,
layer1_node21_MUX_bit_math_h_l959_c3_0003_return_output);

-- layer1_node22_MUX_bit_math_h_l970_c3_fb2c
layer1_node22_MUX_bit_math_h_l970_c3_fb2c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node22_MUX_bit_math_h_l970_c3_fb2c_cond,
layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iftrue,
layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iffalse,
layer1_node22_MUX_bit_math_h_l970_c3_fb2c_return_output);

-- layer1_node23_MUX_bit_math_h_l981_c3_c1f3
layer1_node23_MUX_bit_math_h_l981_c3_c1f3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node23_MUX_bit_math_h_l981_c3_c1f3_cond,
layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iftrue,
layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iffalse,
layer1_node23_MUX_bit_math_h_l981_c3_c1f3_return_output);

-- layer1_node24_MUX_bit_math_h_l992_c3_1884
layer1_node24_MUX_bit_math_h_l992_c3_1884 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node24_MUX_bit_math_h_l992_c3_1884_cond,
layer1_node24_MUX_bit_math_h_l992_c3_1884_iftrue,
layer1_node24_MUX_bit_math_h_l992_c3_1884_iffalse,
layer1_node24_MUX_bit_math_h_l992_c3_1884_return_output);

-- layer1_node25_MUX_bit_math_h_l1003_c3_371a
layer1_node25_MUX_bit_math_h_l1003_c3_371a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node25_MUX_bit_math_h_l1003_c3_371a_cond,
layer1_node25_MUX_bit_math_h_l1003_c3_371a_iftrue,
layer1_node25_MUX_bit_math_h_l1003_c3_371a_iffalse,
layer1_node25_MUX_bit_math_h_l1003_c3_371a_return_output);

-- layer1_node26_MUX_bit_math_h_l1014_c3_b858
layer1_node26_MUX_bit_math_h_l1014_c3_b858 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node26_MUX_bit_math_h_l1014_c3_b858_cond,
layer1_node26_MUX_bit_math_h_l1014_c3_b858_iftrue,
layer1_node26_MUX_bit_math_h_l1014_c3_b858_iffalse,
layer1_node26_MUX_bit_math_h_l1014_c3_b858_return_output);

-- layer1_node27_MUX_bit_math_h_l1025_c3_d07c
layer1_node27_MUX_bit_math_h_l1025_c3_d07c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node27_MUX_bit_math_h_l1025_c3_d07c_cond,
layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iftrue,
layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iffalse,
layer1_node27_MUX_bit_math_h_l1025_c3_d07c_return_output);

-- layer1_node28_MUX_bit_math_h_l1036_c3_d560
layer1_node28_MUX_bit_math_h_l1036_c3_d560 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node28_MUX_bit_math_h_l1036_c3_d560_cond,
layer1_node28_MUX_bit_math_h_l1036_c3_d560_iftrue,
layer1_node28_MUX_bit_math_h_l1036_c3_d560_iffalse,
layer1_node28_MUX_bit_math_h_l1036_c3_d560_return_output);

-- layer1_node29_MUX_bit_math_h_l1047_c3_9f00
layer1_node29_MUX_bit_math_h_l1047_c3_9f00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node29_MUX_bit_math_h_l1047_c3_9f00_cond,
layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iftrue,
layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iffalse,
layer1_node29_MUX_bit_math_h_l1047_c3_9f00_return_output);

-- layer1_node30_MUX_bit_math_h_l1058_c3_e6cc
layer1_node30_MUX_bit_math_h_l1058_c3_e6cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_cond,
layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iftrue,
layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iffalse,
layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_return_output);

-- layer1_node31_MUX_bit_math_h_l1069_c3_b1c7
layer1_node31_MUX_bit_math_h_l1069_c3_b1c7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_cond,
layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iftrue,
layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iffalse,
layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_return_output);

-- layer2_node0_MUX_bit_math_h_l1086_c3_f3d3
layer2_node0_MUX_bit_math_h_l1086_c3_f3d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_cond,
layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iftrue,
layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iffalse,
layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_return_output);

-- layer2_node1_MUX_bit_math_h_l1097_c3_7335
layer2_node1_MUX_bit_math_h_l1097_c3_7335 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l1097_c3_7335_cond,
layer2_node1_MUX_bit_math_h_l1097_c3_7335_iftrue,
layer2_node1_MUX_bit_math_h_l1097_c3_7335_iffalse,
layer2_node1_MUX_bit_math_h_l1097_c3_7335_return_output);

-- layer2_node2_MUX_bit_math_h_l1108_c3_bb5a
layer2_node2_MUX_bit_math_h_l1108_c3_bb5a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_cond,
layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iftrue,
layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iffalse,
layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_return_output);

-- layer2_node3_MUX_bit_math_h_l1119_c3_95be
layer2_node3_MUX_bit_math_h_l1119_c3_95be : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node3_MUX_bit_math_h_l1119_c3_95be_cond,
layer2_node3_MUX_bit_math_h_l1119_c3_95be_iftrue,
layer2_node3_MUX_bit_math_h_l1119_c3_95be_iffalse,
layer2_node3_MUX_bit_math_h_l1119_c3_95be_return_output);

-- layer2_node4_MUX_bit_math_h_l1130_c3_0608
layer2_node4_MUX_bit_math_h_l1130_c3_0608 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node4_MUX_bit_math_h_l1130_c3_0608_cond,
layer2_node4_MUX_bit_math_h_l1130_c3_0608_iftrue,
layer2_node4_MUX_bit_math_h_l1130_c3_0608_iffalse,
layer2_node4_MUX_bit_math_h_l1130_c3_0608_return_output);

-- layer2_node5_MUX_bit_math_h_l1141_c3_a965
layer2_node5_MUX_bit_math_h_l1141_c3_a965 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node5_MUX_bit_math_h_l1141_c3_a965_cond,
layer2_node5_MUX_bit_math_h_l1141_c3_a965_iftrue,
layer2_node5_MUX_bit_math_h_l1141_c3_a965_iffalse,
layer2_node5_MUX_bit_math_h_l1141_c3_a965_return_output);

-- layer2_node6_MUX_bit_math_h_l1152_c3_be4a
layer2_node6_MUX_bit_math_h_l1152_c3_be4a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node6_MUX_bit_math_h_l1152_c3_be4a_cond,
layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iftrue,
layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iffalse,
layer2_node6_MUX_bit_math_h_l1152_c3_be4a_return_output);

-- layer2_node7_MUX_bit_math_h_l1163_c3_4bab
layer2_node7_MUX_bit_math_h_l1163_c3_4bab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node7_MUX_bit_math_h_l1163_c3_4bab_cond,
layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iftrue,
layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iffalse,
layer2_node7_MUX_bit_math_h_l1163_c3_4bab_return_output);

-- layer2_node8_MUX_bit_math_h_l1174_c3_24ff
layer2_node8_MUX_bit_math_h_l1174_c3_24ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node8_MUX_bit_math_h_l1174_c3_24ff_cond,
layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iftrue,
layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iffalse,
layer2_node8_MUX_bit_math_h_l1174_c3_24ff_return_output);

-- layer2_node9_MUX_bit_math_h_l1185_c3_e581
layer2_node9_MUX_bit_math_h_l1185_c3_e581 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node9_MUX_bit_math_h_l1185_c3_e581_cond,
layer2_node9_MUX_bit_math_h_l1185_c3_e581_iftrue,
layer2_node9_MUX_bit_math_h_l1185_c3_e581_iffalse,
layer2_node9_MUX_bit_math_h_l1185_c3_e581_return_output);

-- layer2_node10_MUX_bit_math_h_l1196_c3_c187
layer2_node10_MUX_bit_math_h_l1196_c3_c187 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node10_MUX_bit_math_h_l1196_c3_c187_cond,
layer2_node10_MUX_bit_math_h_l1196_c3_c187_iftrue,
layer2_node10_MUX_bit_math_h_l1196_c3_c187_iffalse,
layer2_node10_MUX_bit_math_h_l1196_c3_c187_return_output);

-- layer2_node11_MUX_bit_math_h_l1207_c3_bafc
layer2_node11_MUX_bit_math_h_l1207_c3_bafc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node11_MUX_bit_math_h_l1207_c3_bafc_cond,
layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iftrue,
layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iffalse,
layer2_node11_MUX_bit_math_h_l1207_c3_bafc_return_output);

-- layer2_node12_MUX_bit_math_h_l1218_c3_c26f
layer2_node12_MUX_bit_math_h_l1218_c3_c26f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node12_MUX_bit_math_h_l1218_c3_c26f_cond,
layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iftrue,
layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iffalse,
layer2_node12_MUX_bit_math_h_l1218_c3_c26f_return_output);

-- layer2_node13_MUX_bit_math_h_l1229_c3_bcb9
layer2_node13_MUX_bit_math_h_l1229_c3_bcb9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_cond,
layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iftrue,
layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iffalse,
layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_return_output);

-- layer2_node14_MUX_bit_math_h_l1240_c3_7be3
layer2_node14_MUX_bit_math_h_l1240_c3_7be3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node14_MUX_bit_math_h_l1240_c3_7be3_cond,
layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iftrue,
layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iffalse,
layer2_node14_MUX_bit_math_h_l1240_c3_7be3_return_output);

-- layer2_node15_MUX_bit_math_h_l1251_c3_1e63
layer2_node15_MUX_bit_math_h_l1251_c3_1e63 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node15_MUX_bit_math_h_l1251_c3_1e63_cond,
layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iftrue,
layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iffalse,
layer2_node15_MUX_bit_math_h_l1251_c3_1e63_return_output);

-- layer3_node0_MUX_bit_math_h_l1268_c3_e356
layer3_node0_MUX_bit_math_h_l1268_c3_e356 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l1268_c3_e356_cond,
layer3_node0_MUX_bit_math_h_l1268_c3_e356_iftrue,
layer3_node0_MUX_bit_math_h_l1268_c3_e356_iffalse,
layer3_node0_MUX_bit_math_h_l1268_c3_e356_return_output);

-- layer3_node1_MUX_bit_math_h_l1279_c3_3873
layer3_node1_MUX_bit_math_h_l1279_c3_3873 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node1_MUX_bit_math_h_l1279_c3_3873_cond,
layer3_node1_MUX_bit_math_h_l1279_c3_3873_iftrue,
layer3_node1_MUX_bit_math_h_l1279_c3_3873_iffalse,
layer3_node1_MUX_bit_math_h_l1279_c3_3873_return_output);

-- layer3_node2_MUX_bit_math_h_l1290_c3_4ec7
layer3_node2_MUX_bit_math_h_l1290_c3_4ec7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_cond,
layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iftrue,
layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iffalse,
layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_return_output);

-- layer3_node3_MUX_bit_math_h_l1301_c3_29f9
layer3_node3_MUX_bit_math_h_l1301_c3_29f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node3_MUX_bit_math_h_l1301_c3_29f9_cond,
layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iftrue,
layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iffalse,
layer3_node3_MUX_bit_math_h_l1301_c3_29f9_return_output);

-- layer3_node4_MUX_bit_math_h_l1312_c3_b484
layer3_node4_MUX_bit_math_h_l1312_c3_b484 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node4_MUX_bit_math_h_l1312_c3_b484_cond,
layer3_node4_MUX_bit_math_h_l1312_c3_b484_iftrue,
layer3_node4_MUX_bit_math_h_l1312_c3_b484_iffalse,
layer3_node4_MUX_bit_math_h_l1312_c3_b484_return_output);

-- layer3_node5_MUX_bit_math_h_l1323_c3_e63b
layer3_node5_MUX_bit_math_h_l1323_c3_e63b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node5_MUX_bit_math_h_l1323_c3_e63b_cond,
layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iftrue,
layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iffalse,
layer3_node5_MUX_bit_math_h_l1323_c3_e63b_return_output);

-- layer3_node6_MUX_bit_math_h_l1334_c3_5def
layer3_node6_MUX_bit_math_h_l1334_c3_5def : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node6_MUX_bit_math_h_l1334_c3_5def_cond,
layer3_node6_MUX_bit_math_h_l1334_c3_5def_iftrue,
layer3_node6_MUX_bit_math_h_l1334_c3_5def_iffalse,
layer3_node6_MUX_bit_math_h_l1334_c3_5def_return_output);

-- layer3_node7_MUX_bit_math_h_l1345_c3_3cb2
layer3_node7_MUX_bit_math_h_l1345_c3_3cb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_cond,
layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iftrue,
layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iffalse,
layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_return_output);

-- layer4_node0_MUX_bit_math_h_l1362_c3_fa41
layer4_node0_MUX_bit_math_h_l1362_c3_fa41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node0_MUX_bit_math_h_l1362_c3_fa41_cond,
layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iftrue,
layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iffalse,
layer4_node0_MUX_bit_math_h_l1362_c3_fa41_return_output);

-- layer4_node1_MUX_bit_math_h_l1373_c3_223f
layer4_node1_MUX_bit_math_h_l1373_c3_223f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node1_MUX_bit_math_h_l1373_c3_223f_cond,
layer4_node1_MUX_bit_math_h_l1373_c3_223f_iftrue,
layer4_node1_MUX_bit_math_h_l1373_c3_223f_iffalse,
layer4_node1_MUX_bit_math_h_l1373_c3_223f_return_output);

-- layer4_node2_MUX_bit_math_h_l1384_c3_470b
layer4_node2_MUX_bit_math_h_l1384_c3_470b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node2_MUX_bit_math_h_l1384_c3_470b_cond,
layer4_node2_MUX_bit_math_h_l1384_c3_470b_iftrue,
layer4_node2_MUX_bit_math_h_l1384_c3_470b_iffalse,
layer4_node2_MUX_bit_math_h_l1384_c3_470b_return_output);

-- layer4_node3_MUX_bit_math_h_l1395_c3_68f4
layer4_node3_MUX_bit_math_h_l1395_c3_68f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node3_MUX_bit_math_h_l1395_c3_68f4_cond,
layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iftrue,
layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iffalse,
layer4_node3_MUX_bit_math_h_l1395_c3_68f4_return_output);

-- layer5_node0_MUX_bit_math_h_l1412_c3_e3bb
layer5_node0_MUX_bit_math_h_l1412_c3_e3bb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_cond,
layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iftrue,
layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iffalse,
layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_return_output);

-- layer5_node1_MUX_bit_math_h_l1423_c3_47e8
layer5_node1_MUX_bit_math_h_l1423_c3_47e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node1_MUX_bit_math_h_l1423_c3_47e8_cond,
layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iftrue,
layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iffalse,
layer5_node1_MUX_bit_math_h_l1423_c3_47e8_return_output);

-- layer6_node0_MUX_bit_math_h_l1440_c3_7682
layer6_node0_MUX_bit_math_h_l1440_c3_7682 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer6_node0_MUX_bit_math_h_l1440_c3_7682_cond,
layer6_node0_MUX_bit_math_h_l1440_c3_7682_iftrue,
layer6_node0_MUX_bit_math_h_l1440_c3_7682_iffalse,
layer6_node0_MUX_bit_math_h_l1440_c3_7682_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 in16,
 in17,
 in18,
 in19,
 in20,
 in21,
 in22,
 in23,
 in24,
 in25,
 in26,
 in27,
 in28,
 in29,
 in30,
 in31,
 in32,
 in33,
 in34,
 in35,
 in36,
 in37,
 in38,
 in39,
 in40,
 in41,
 in42,
 in43,
 in44,
 in45,
 in46,
 in47,
 in48,
 in49,
 in50,
 in51,
 in52,
 in53,
 in54,
 in55,
 in56,
 in57,
 in58,
 in59,
 in60,
 in61,
 in62,
 in63,
 in64,
 in65,
 in66,
 in67,
 in68,
 in69,
 in70,
 in71,
 in72,
 in73,
 in74,
 in75,
 in76,
 in77,
 in78,
 in79,
 in80,
 in81,
 in82,
 in83,
 in84,
 in85,
 in86,
 in87,
 in88,
 in89,
 in90,
 in91,
 in92,
 in93,
 in94,
 in95,
 in96,
 in97,
 in98,
 in99,
 in100,
 in101,
 in102,
 in103,
 in104,
 in105,
 in106,
 in107,
 in108,
 in109,
 in110,
 in111,
 in112,
 in113,
 in114,
 in115,
 in116,
 in117,
 in118,
 in119,
 in120,
 in121,
 in122,
 in123,
 in124,
 in125,
 in126,
 in127,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_70c7_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_dc12_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_3404_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_cc01_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_7793_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_2acd_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_494b_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_daab_return_output,
 layer0_node8_MUX_bit_math_h_l106_c3_d50d_return_output,
 layer0_node9_MUX_bit_math_h_l117_c3_c9ee_return_output,
 layer0_node10_MUX_bit_math_h_l128_c3_06d1_return_output,
 layer0_node11_MUX_bit_math_h_l139_c3_13dc_return_output,
 layer0_node12_MUX_bit_math_h_l150_c3_af2c_return_output,
 layer0_node13_MUX_bit_math_h_l161_c3_c865_return_output,
 layer0_node14_MUX_bit_math_h_l172_c3_1937_return_output,
 layer0_node15_MUX_bit_math_h_l183_c3_6211_return_output,
 layer0_node16_MUX_bit_math_h_l194_c3_6e24_return_output,
 layer0_node17_MUX_bit_math_h_l205_c3_4b2c_return_output,
 layer0_node18_MUX_bit_math_h_l216_c3_0b83_return_output,
 layer0_node19_MUX_bit_math_h_l227_c3_1e36_return_output,
 layer0_node20_MUX_bit_math_h_l238_c3_5458_return_output,
 layer0_node21_MUX_bit_math_h_l249_c3_c173_return_output,
 layer0_node22_MUX_bit_math_h_l260_c3_fce5_return_output,
 layer0_node23_MUX_bit_math_h_l271_c3_a82d_return_output,
 layer0_node24_MUX_bit_math_h_l282_c3_6611_return_output,
 layer0_node25_MUX_bit_math_h_l293_c3_b4b9_return_output,
 layer0_node26_MUX_bit_math_h_l304_c3_2bce_return_output,
 layer0_node27_MUX_bit_math_h_l315_c3_7789_return_output,
 layer0_node28_MUX_bit_math_h_l326_c3_098d_return_output,
 layer0_node29_MUX_bit_math_h_l337_c3_9c87_return_output,
 layer0_node30_MUX_bit_math_h_l348_c3_6b0d_return_output,
 layer0_node31_MUX_bit_math_h_l359_c3_5065_return_output,
 layer0_node32_MUX_bit_math_h_l370_c3_4893_return_output,
 layer0_node33_MUX_bit_math_h_l381_c3_8132_return_output,
 layer0_node34_MUX_bit_math_h_l392_c3_59bd_return_output,
 layer0_node35_MUX_bit_math_h_l403_c3_6326_return_output,
 layer0_node36_MUX_bit_math_h_l414_c3_7348_return_output,
 layer0_node37_MUX_bit_math_h_l425_c3_f929_return_output,
 layer0_node38_MUX_bit_math_h_l436_c3_d3a0_return_output,
 layer0_node39_MUX_bit_math_h_l447_c3_7b35_return_output,
 layer0_node40_MUX_bit_math_h_l458_c3_426b_return_output,
 layer0_node41_MUX_bit_math_h_l469_c3_47d5_return_output,
 layer0_node42_MUX_bit_math_h_l480_c3_50c3_return_output,
 layer0_node43_MUX_bit_math_h_l491_c3_6ed7_return_output,
 layer0_node44_MUX_bit_math_h_l502_c3_84a4_return_output,
 layer0_node45_MUX_bit_math_h_l513_c3_552e_return_output,
 layer0_node46_MUX_bit_math_h_l524_c3_42cd_return_output,
 layer0_node47_MUX_bit_math_h_l535_c3_18b2_return_output,
 layer0_node48_MUX_bit_math_h_l546_c3_e9fe_return_output,
 layer0_node49_MUX_bit_math_h_l557_c3_68c1_return_output,
 layer0_node50_MUX_bit_math_h_l568_c3_8ec7_return_output,
 layer0_node51_MUX_bit_math_h_l579_c3_5985_return_output,
 layer0_node52_MUX_bit_math_h_l590_c3_90c2_return_output,
 layer0_node53_MUX_bit_math_h_l601_c3_5a9e_return_output,
 layer0_node54_MUX_bit_math_h_l612_c3_235a_return_output,
 layer0_node55_MUX_bit_math_h_l623_c3_1dea_return_output,
 layer0_node56_MUX_bit_math_h_l634_c3_f6e3_return_output,
 layer0_node57_MUX_bit_math_h_l645_c3_eeb0_return_output,
 layer0_node58_MUX_bit_math_h_l656_c3_b995_return_output,
 layer0_node59_MUX_bit_math_h_l667_c3_b104_return_output,
 layer0_node60_MUX_bit_math_h_l678_c3_7571_return_output,
 layer0_node61_MUX_bit_math_h_l689_c3_580e_return_output,
 layer0_node62_MUX_bit_math_h_l700_c3_9f5f_return_output,
 layer0_node63_MUX_bit_math_h_l711_c3_17f2_return_output,
 layer1_node0_MUX_bit_math_h_l728_c3_23e3_return_output,
 layer1_node1_MUX_bit_math_h_l739_c3_57f6_return_output,
 layer1_node2_MUX_bit_math_h_l750_c3_b86b_return_output,
 layer1_node3_MUX_bit_math_h_l761_c3_2586_return_output,
 layer1_node4_MUX_bit_math_h_l772_c3_857f_return_output,
 layer1_node5_MUX_bit_math_h_l783_c3_f8bc_return_output,
 layer1_node6_MUX_bit_math_h_l794_c3_f4dd_return_output,
 layer1_node7_MUX_bit_math_h_l805_c3_e535_return_output,
 layer1_node8_MUX_bit_math_h_l816_c3_e51d_return_output,
 layer1_node9_MUX_bit_math_h_l827_c3_4f17_return_output,
 layer1_node10_MUX_bit_math_h_l838_c3_8caa_return_output,
 layer1_node11_MUX_bit_math_h_l849_c3_c418_return_output,
 layer1_node12_MUX_bit_math_h_l860_c3_3ea5_return_output,
 layer1_node13_MUX_bit_math_h_l871_c3_66e4_return_output,
 layer1_node14_MUX_bit_math_h_l882_c3_5e4a_return_output,
 layer1_node15_MUX_bit_math_h_l893_c3_faee_return_output,
 layer1_node16_MUX_bit_math_h_l904_c3_1e1f_return_output,
 layer1_node17_MUX_bit_math_h_l915_c3_bbc7_return_output,
 layer1_node18_MUX_bit_math_h_l926_c3_15bb_return_output,
 layer1_node19_MUX_bit_math_h_l937_c3_3ad6_return_output,
 layer1_node20_MUX_bit_math_h_l948_c3_d497_return_output,
 layer1_node21_MUX_bit_math_h_l959_c3_0003_return_output,
 layer1_node22_MUX_bit_math_h_l970_c3_fb2c_return_output,
 layer1_node23_MUX_bit_math_h_l981_c3_c1f3_return_output,
 layer1_node24_MUX_bit_math_h_l992_c3_1884_return_output,
 layer1_node25_MUX_bit_math_h_l1003_c3_371a_return_output,
 layer1_node26_MUX_bit_math_h_l1014_c3_b858_return_output,
 layer1_node27_MUX_bit_math_h_l1025_c3_d07c_return_output,
 layer1_node28_MUX_bit_math_h_l1036_c3_d560_return_output,
 layer1_node29_MUX_bit_math_h_l1047_c3_9f00_return_output,
 layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_return_output,
 layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_return_output,
 layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_return_output,
 layer2_node1_MUX_bit_math_h_l1097_c3_7335_return_output,
 layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_return_output,
 layer2_node3_MUX_bit_math_h_l1119_c3_95be_return_output,
 layer2_node4_MUX_bit_math_h_l1130_c3_0608_return_output,
 layer2_node5_MUX_bit_math_h_l1141_c3_a965_return_output,
 layer2_node6_MUX_bit_math_h_l1152_c3_be4a_return_output,
 layer2_node7_MUX_bit_math_h_l1163_c3_4bab_return_output,
 layer2_node8_MUX_bit_math_h_l1174_c3_24ff_return_output,
 layer2_node9_MUX_bit_math_h_l1185_c3_e581_return_output,
 layer2_node10_MUX_bit_math_h_l1196_c3_c187_return_output,
 layer2_node11_MUX_bit_math_h_l1207_c3_bafc_return_output,
 layer2_node12_MUX_bit_math_h_l1218_c3_c26f_return_output,
 layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_return_output,
 layer2_node14_MUX_bit_math_h_l1240_c3_7be3_return_output,
 layer2_node15_MUX_bit_math_h_l1251_c3_1e63_return_output,
 layer3_node0_MUX_bit_math_h_l1268_c3_e356_return_output,
 layer3_node1_MUX_bit_math_h_l1279_c3_3873_return_output,
 layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_return_output,
 layer3_node3_MUX_bit_math_h_l1301_c3_29f9_return_output,
 layer3_node4_MUX_bit_math_h_l1312_c3_b484_return_output,
 layer3_node5_MUX_bit_math_h_l1323_c3_e63b_return_output,
 layer3_node6_MUX_bit_math_h_l1334_c3_5def_return_output,
 layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_return_output,
 layer4_node0_MUX_bit_math_h_l1362_c3_fa41_return_output,
 layer4_node1_MUX_bit_math_h_l1373_c3_223f_return_output,
 layer4_node2_MUX_bit_math_h_l1384_c3_470b_return_output,
 layer4_node3_MUX_bit_math_h_l1395_c3_68f4_return_output,
 layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_return_output,
 layer5_node1_MUX_bit_math_h_l1423_c3_47e8_return_output,
 layer6_node0_MUX_bit_math_h_l1440_c3_7682_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(7 downto 0);
 variable VAR_sel : unsigned(6 downto 0);
 variable VAR_in0 : unsigned(7 downto 0);
 variable VAR_in1 : unsigned(7 downto 0);
 variable VAR_in2 : unsigned(7 downto 0);
 variable VAR_in3 : unsigned(7 downto 0);
 variable VAR_in4 : unsigned(7 downto 0);
 variable VAR_in5 : unsigned(7 downto 0);
 variable VAR_in6 : unsigned(7 downto 0);
 variable VAR_in7 : unsigned(7 downto 0);
 variable VAR_in8 : unsigned(7 downto 0);
 variable VAR_in9 : unsigned(7 downto 0);
 variable VAR_in10 : unsigned(7 downto 0);
 variable VAR_in11 : unsigned(7 downto 0);
 variable VAR_in12 : unsigned(7 downto 0);
 variable VAR_in13 : unsigned(7 downto 0);
 variable VAR_in14 : unsigned(7 downto 0);
 variable VAR_in15 : unsigned(7 downto 0);
 variable VAR_in16 : unsigned(7 downto 0);
 variable VAR_in17 : unsigned(7 downto 0);
 variable VAR_in18 : unsigned(7 downto 0);
 variable VAR_in19 : unsigned(7 downto 0);
 variable VAR_in20 : unsigned(7 downto 0);
 variable VAR_in21 : unsigned(7 downto 0);
 variable VAR_in22 : unsigned(7 downto 0);
 variable VAR_in23 : unsigned(7 downto 0);
 variable VAR_in24 : unsigned(7 downto 0);
 variable VAR_in25 : unsigned(7 downto 0);
 variable VAR_in26 : unsigned(7 downto 0);
 variable VAR_in27 : unsigned(7 downto 0);
 variable VAR_in28 : unsigned(7 downto 0);
 variable VAR_in29 : unsigned(7 downto 0);
 variable VAR_in30 : unsigned(7 downto 0);
 variable VAR_in31 : unsigned(7 downto 0);
 variable VAR_in32 : unsigned(7 downto 0);
 variable VAR_in33 : unsigned(7 downto 0);
 variable VAR_in34 : unsigned(7 downto 0);
 variable VAR_in35 : unsigned(7 downto 0);
 variable VAR_in36 : unsigned(7 downto 0);
 variable VAR_in37 : unsigned(7 downto 0);
 variable VAR_in38 : unsigned(7 downto 0);
 variable VAR_in39 : unsigned(7 downto 0);
 variable VAR_in40 : unsigned(7 downto 0);
 variable VAR_in41 : unsigned(7 downto 0);
 variable VAR_in42 : unsigned(7 downto 0);
 variable VAR_in43 : unsigned(7 downto 0);
 variable VAR_in44 : unsigned(7 downto 0);
 variable VAR_in45 : unsigned(7 downto 0);
 variable VAR_in46 : unsigned(7 downto 0);
 variable VAR_in47 : unsigned(7 downto 0);
 variable VAR_in48 : unsigned(7 downto 0);
 variable VAR_in49 : unsigned(7 downto 0);
 variable VAR_in50 : unsigned(7 downto 0);
 variable VAR_in51 : unsigned(7 downto 0);
 variable VAR_in52 : unsigned(7 downto 0);
 variable VAR_in53 : unsigned(7 downto 0);
 variable VAR_in54 : unsigned(7 downto 0);
 variable VAR_in55 : unsigned(7 downto 0);
 variable VAR_in56 : unsigned(7 downto 0);
 variable VAR_in57 : unsigned(7 downto 0);
 variable VAR_in58 : unsigned(7 downto 0);
 variable VAR_in59 : unsigned(7 downto 0);
 variable VAR_in60 : unsigned(7 downto 0);
 variable VAR_in61 : unsigned(7 downto 0);
 variable VAR_in62 : unsigned(7 downto 0);
 variable VAR_in63 : unsigned(7 downto 0);
 variable VAR_in64 : unsigned(7 downto 0);
 variable VAR_in65 : unsigned(7 downto 0);
 variable VAR_in66 : unsigned(7 downto 0);
 variable VAR_in67 : unsigned(7 downto 0);
 variable VAR_in68 : unsigned(7 downto 0);
 variable VAR_in69 : unsigned(7 downto 0);
 variable VAR_in70 : unsigned(7 downto 0);
 variable VAR_in71 : unsigned(7 downto 0);
 variable VAR_in72 : unsigned(7 downto 0);
 variable VAR_in73 : unsigned(7 downto 0);
 variable VAR_in74 : unsigned(7 downto 0);
 variable VAR_in75 : unsigned(7 downto 0);
 variable VAR_in76 : unsigned(7 downto 0);
 variable VAR_in77 : unsigned(7 downto 0);
 variable VAR_in78 : unsigned(7 downto 0);
 variable VAR_in79 : unsigned(7 downto 0);
 variable VAR_in80 : unsigned(7 downto 0);
 variable VAR_in81 : unsigned(7 downto 0);
 variable VAR_in82 : unsigned(7 downto 0);
 variable VAR_in83 : unsigned(7 downto 0);
 variable VAR_in84 : unsigned(7 downto 0);
 variable VAR_in85 : unsigned(7 downto 0);
 variable VAR_in86 : unsigned(7 downto 0);
 variable VAR_in87 : unsigned(7 downto 0);
 variable VAR_in88 : unsigned(7 downto 0);
 variable VAR_in89 : unsigned(7 downto 0);
 variable VAR_in90 : unsigned(7 downto 0);
 variable VAR_in91 : unsigned(7 downto 0);
 variable VAR_in92 : unsigned(7 downto 0);
 variable VAR_in93 : unsigned(7 downto 0);
 variable VAR_in94 : unsigned(7 downto 0);
 variable VAR_in95 : unsigned(7 downto 0);
 variable VAR_in96 : unsigned(7 downto 0);
 variable VAR_in97 : unsigned(7 downto 0);
 variable VAR_in98 : unsigned(7 downto 0);
 variable VAR_in99 : unsigned(7 downto 0);
 variable VAR_in100 : unsigned(7 downto 0);
 variable VAR_in101 : unsigned(7 downto 0);
 variable VAR_in102 : unsigned(7 downto 0);
 variable VAR_in103 : unsigned(7 downto 0);
 variable VAR_in104 : unsigned(7 downto 0);
 variable VAR_in105 : unsigned(7 downto 0);
 variable VAR_in106 : unsigned(7 downto 0);
 variable VAR_in107 : unsigned(7 downto 0);
 variable VAR_in108 : unsigned(7 downto 0);
 variable VAR_in109 : unsigned(7 downto 0);
 variable VAR_in110 : unsigned(7 downto 0);
 variable VAR_in111 : unsigned(7 downto 0);
 variable VAR_in112 : unsigned(7 downto 0);
 variable VAR_in113 : unsigned(7 downto 0);
 variable VAR_in114 : unsigned(7 downto 0);
 variable VAR_in115 : unsigned(7 downto 0);
 variable VAR_in116 : unsigned(7 downto 0);
 variable VAR_in117 : unsigned(7 downto 0);
 variable VAR_in118 : unsigned(7 downto 0);
 variable VAR_in119 : unsigned(7 downto 0);
 variable VAR_in120 : unsigned(7 downto 0);
 variable VAR_in121 : unsigned(7 downto 0);
 variable VAR_in122 : unsigned(7 downto 0);
 variable VAR_in123 : unsigned(7 downto 0);
 variable VAR_in124 : unsigned(7 downto 0);
 variable VAR_in125 : unsigned(7 downto 0);
 variable VAR_in126 : unsigned(7 downto 0);
 variable VAR_in127 : unsigned(7 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_cond : unsigned(0 downto 0);
 variable VAR_layer0_node8 : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node9 : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_cond : unsigned(0 downto 0);
 variable VAR_layer0_node10 : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node11 : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_cond : unsigned(0 downto 0);
 variable VAR_layer0_node12 : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node13 : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_cond : unsigned(0 downto 0);
 variable VAR_layer0_node14 : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_cond : unsigned(0 downto 0);
 variable VAR_layer0_node15 : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_cond : unsigned(0 downto 0);
 variable VAR_layer0_node16 : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_cond : unsigned(0 downto 0);
 variable VAR_layer0_node17 : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node18 : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_cond : unsigned(0 downto 0);
 variable VAR_layer0_node19 : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_cond : unsigned(0 downto 0);
 variable VAR_layer0_node20 : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_cond : unsigned(0 downto 0);
 variable VAR_layer0_node21 : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_cond : unsigned(0 downto 0);
 variable VAR_layer0_node22 : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_cond : unsigned(0 downto 0);
 variable VAR_layer0_node23 : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node24 : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_cond : unsigned(0 downto 0);
 variable VAR_layer0_node25 : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node26 : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_cond : unsigned(0 downto 0);
 variable VAR_layer0_node27 : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_cond : unsigned(0 downto 0);
 variable VAR_layer0_node28 : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node29 : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_cond : unsigned(0 downto 0);
 variable VAR_layer0_node30 : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node31 : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_cond : unsigned(0 downto 0);
 variable VAR_layer0_node32 : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_cond : unsigned(0 downto 0);
 variable VAR_layer0_node33 : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_cond : unsigned(0 downto 0);
 variable VAR_layer0_node34 : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_cond : unsigned(0 downto 0);
 variable VAR_layer0_node35 : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_cond : unsigned(0 downto 0);
 variable VAR_layer0_node36 : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_cond : unsigned(0 downto 0);
 variable VAR_layer0_node37 : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_cond : unsigned(0 downto 0);
 variable VAR_layer0_node38 : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_cond : unsigned(0 downto 0);
 variable VAR_layer0_node39 : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_cond : unsigned(0 downto 0);
 variable VAR_layer0_node40 : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node41 : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_cond : unsigned(0 downto 0);
 variable VAR_layer0_node42 : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node43 : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node44 : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_cond : unsigned(0 downto 0);
 variable VAR_layer0_node45 : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node46 : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_cond : unsigned(0 downto 0);
 variable VAR_layer0_node47 : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node48 : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_cond : unsigned(0 downto 0);
 variable VAR_layer0_node49 : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node50 : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node51 : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_cond : unsigned(0 downto 0);
 variable VAR_layer0_node52 : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node53 : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node54 : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node55 : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_cond : unsigned(0 downto 0);
 variable VAR_layer0_node56 : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node57 : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_cond : unsigned(0 downto 0);
 variable VAR_layer0_node58 : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_cond : unsigned(0 downto 0);
 variable VAR_layer0_node59 : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_cond : unsigned(0 downto 0);
 variable VAR_layer0_node60 : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_cond : unsigned(0 downto 0);
 variable VAR_layer0_node61 : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node62 : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_cond : unsigned(0 downto 0);
 variable VAR_layer0_node63 : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_cond : unsigned(0 downto 0);
 variable VAR_layer1_node4 : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node5 : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_cond : unsigned(0 downto 0);
 variable VAR_layer1_node6 : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_cond : unsigned(0 downto 0);
 variable VAR_layer1_node7 : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_cond : unsigned(0 downto 0);
 variable VAR_layer1_node8 : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_cond : unsigned(0 downto 0);
 variable VAR_layer1_node9 : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_cond : unsigned(0 downto 0);
 variable VAR_layer1_node10 : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_cond : unsigned(0 downto 0);
 variable VAR_layer1_node11 : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_cond : unsigned(0 downto 0);
 variable VAR_layer1_node12 : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_cond : unsigned(0 downto 0);
 variable VAR_layer1_node13 : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_cond : unsigned(0 downto 0);
 variable VAR_layer1_node14 : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_cond : unsigned(0 downto 0);
 variable VAR_layer1_node15 : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_cond : unsigned(0 downto 0);
 variable VAR_layer1_node16 : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node17 : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_cond : unsigned(0 downto 0);
 variable VAR_layer1_node18 : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_cond : unsigned(0 downto 0);
 variable VAR_layer1_node19 : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_cond : unsigned(0 downto 0);
 variable VAR_layer1_node20 : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_cond : unsigned(0 downto 0);
 variable VAR_layer1_node21 : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_cond : unsigned(0 downto 0);
 variable VAR_layer1_node22 : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_cond : unsigned(0 downto 0);
 variable VAR_layer1_node23 : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_cond : unsigned(0 downto 0);
 variable VAR_layer1_node24 : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_cond : unsigned(0 downto 0);
 variable VAR_layer1_node25 : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_cond : unsigned(0 downto 0);
 variable VAR_layer1_node26 : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_cond : unsigned(0 downto 0);
 variable VAR_layer1_node27 : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_cond : unsigned(0 downto 0);
 variable VAR_layer1_node28 : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_cond : unsigned(0 downto 0);
 variable VAR_layer1_node29 : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_cond : unsigned(0 downto 0);
 variable VAR_layer1_node30 : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_cond : unsigned(0 downto 0);
 variable VAR_layer1_node31 : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_cond : unsigned(0 downto 0);
 variable VAR_layer2_node2 : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_cond : unsigned(0 downto 0);
 variable VAR_layer2_node3 : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_cond : unsigned(0 downto 0);
 variable VAR_layer2_node4 : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_cond : unsigned(0 downto 0);
 variable VAR_layer2_node5 : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_cond : unsigned(0 downto 0);
 variable VAR_layer2_node6 : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_cond : unsigned(0 downto 0);
 variable VAR_layer2_node7 : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_cond : unsigned(0 downto 0);
 variable VAR_layer2_node8 : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_cond : unsigned(0 downto 0);
 variable VAR_layer2_node9 : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_cond : unsigned(0 downto 0);
 variable VAR_layer2_node10 : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_cond : unsigned(0 downto 0);
 variable VAR_layer2_node11 : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_cond : unsigned(0 downto 0);
 variable VAR_layer2_node12 : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_cond : unsigned(0 downto 0);
 variable VAR_layer2_node13 : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_cond : unsigned(0 downto 0);
 variable VAR_layer2_node14 : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_cond : unsigned(0 downto 0);
 variable VAR_layer2_node15 : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_cond : unsigned(0 downto 0);
 variable VAR_layer3_node1 : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_cond : unsigned(0 downto 0);
 variable VAR_layer3_node2 : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_cond : unsigned(0 downto 0);
 variable VAR_layer3_node3 : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_cond : unsigned(0 downto 0);
 variable VAR_layer3_node4 : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_cond : unsigned(0 downto 0);
 variable VAR_layer3_node5 : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_cond : unsigned(0 downto 0);
 variable VAR_layer3_node6 : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_cond : unsigned(0 downto 0);
 variable VAR_layer3_node7 : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_cond : unsigned(0 downto 0);
 variable VAR_sel4 : unsigned(0 downto 0);
 variable VAR_uint7_4_4_bit_math_h_l1358_c10_7de3_return_output : unsigned(0 downto 0);
 variable VAR_layer4_node0 : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_cond : unsigned(0 downto 0);
 variable VAR_layer4_node1 : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_cond : unsigned(0 downto 0);
 variable VAR_layer4_node2 : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_cond : unsigned(0 downto 0);
 variable VAR_layer4_node3 : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_cond : unsigned(0 downto 0);
 variable VAR_sel5 : unsigned(0 downto 0);
 variable VAR_uint7_5_5_bit_math_h_l1408_c10_6715_return_output : unsigned(0 downto 0);
 variable VAR_layer5_node0 : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_cond : unsigned(0 downto 0);
 variable VAR_layer5_node1 : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_cond : unsigned(0 downto 0);
 variable VAR_sel6 : unsigned(0 downto 0);
 variable VAR_uint7_6_6_bit_math_h_l1436_c10_2546_return_output : unsigned(0 downto 0);
 variable VAR_layer6_node0 : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_iftrue : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_iffalse : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_return_output : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;
     VAR_in16 := in16;
     VAR_in17 := in17;
     VAR_in18 := in18;
     VAR_in19 := in19;
     VAR_in20 := in20;
     VAR_in21 := in21;
     VAR_in22 := in22;
     VAR_in23 := in23;
     VAR_in24 := in24;
     VAR_in25 := in25;
     VAR_in26 := in26;
     VAR_in27 := in27;
     VAR_in28 := in28;
     VAR_in29 := in29;
     VAR_in30 := in30;
     VAR_in31 := in31;
     VAR_in32 := in32;
     VAR_in33 := in33;
     VAR_in34 := in34;
     VAR_in35 := in35;
     VAR_in36 := in36;
     VAR_in37 := in37;
     VAR_in38 := in38;
     VAR_in39 := in39;
     VAR_in40 := in40;
     VAR_in41 := in41;
     VAR_in42 := in42;
     VAR_in43 := in43;
     VAR_in44 := in44;
     VAR_in45 := in45;
     VAR_in46 := in46;
     VAR_in47 := in47;
     VAR_in48 := in48;
     VAR_in49 := in49;
     VAR_in50 := in50;
     VAR_in51 := in51;
     VAR_in52 := in52;
     VAR_in53 := in53;
     VAR_in54 := in54;
     VAR_in55 := in55;
     VAR_in56 := in56;
     VAR_in57 := in57;
     VAR_in58 := in58;
     VAR_in59 := in59;
     VAR_in60 := in60;
     VAR_in61 := in61;
     VAR_in62 := in62;
     VAR_in63 := in63;
     VAR_in64 := in64;
     VAR_in65 := in65;
     VAR_in66 := in66;
     VAR_in67 := in67;
     VAR_in68 := in68;
     VAR_in69 := in69;
     VAR_in70 := in70;
     VAR_in71 := in71;
     VAR_in72 := in72;
     VAR_in73 := in73;
     VAR_in74 := in74;
     VAR_in75 := in75;
     VAR_in76 := in76;
     VAR_in77 := in77;
     VAR_in78 := in78;
     VAR_in79 := in79;
     VAR_in80 := in80;
     VAR_in81 := in81;
     VAR_in82 := in82;
     VAR_in83 := in83;
     VAR_in84 := in84;
     VAR_in85 := in85;
     VAR_in86 := in86;
     VAR_in87 := in87;
     VAR_in88 := in88;
     VAR_in89 := in89;
     VAR_in90 := in90;
     VAR_in91 := in91;
     VAR_in92 := in92;
     VAR_in93 := in93;
     VAR_in94 := in94;
     VAR_in95 := in95;
     VAR_in96 := in96;
     VAR_in97 := in97;
     VAR_in98 := in98;
     VAR_in99 := in99;
     VAR_in100 := in100;
     VAR_in101 := in101;
     VAR_in102 := in102;
     VAR_in103 := in103;
     VAR_in104 := in104;
     VAR_in105 := in105;
     VAR_in106 := in106;
     VAR_in107 := in107;
     VAR_in108 := in108;
     VAR_in109 := in109;
     VAR_in110 := in110;
     VAR_in111 := in111;
     VAR_in112 := in112;
     VAR_in113 := in113;
     VAR_in114 := in114;
     VAR_in115 := in115;
     VAR_in116 := in116;
     VAR_in117 := in117;
     VAR_in118 := in118;
     VAR_in119 := in119;
     VAR_in120 := in120;
     VAR_in121 := in121;
     VAR_in122 := in122;
     VAR_in123 := in123;
     VAR_in124 := in124;
     VAR_in125 := in125;
     VAR_in126 := in126;
     VAR_in127 := in127;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_iffalse := VAR_in10;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iffalse := VAR_in100;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iftrue := VAR_in101;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_iffalse := VAR_in102;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_iftrue := VAR_in103;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_iffalse := VAR_in104;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_iftrue := VAR_in105;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iffalse := VAR_in106;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iftrue := VAR_in107;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_iffalse := VAR_in108;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_iftrue := VAR_in109;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_iftrue := VAR_in11;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_iffalse := VAR_in110;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_iftrue := VAR_in111;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iffalse := VAR_in112;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iftrue := VAR_in113;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iffalse := VAR_in114;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iftrue := VAR_in115;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_iffalse := VAR_in116;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_iftrue := VAR_in117;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_iffalse := VAR_in118;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_iftrue := VAR_in119;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_iffalse := VAR_in12;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_iffalse := VAR_in120;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_iftrue := VAR_in121;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_iffalse := VAR_in122;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_iftrue := VAR_in123;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iffalse := VAR_in124;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iftrue := VAR_in125;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_iffalse := VAR_in126;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_iftrue := VAR_in127;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_iftrue := VAR_in15;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_iffalse := VAR_in16;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_iftrue := VAR_in17;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iffalse := VAR_in18;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iftrue := VAR_in19;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_iffalse := VAR_in2;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_iffalse := VAR_in20;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_iftrue := VAR_in21;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_iffalse := VAR_in22;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_iftrue := VAR_in23;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_iffalse := VAR_in24;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_iftrue := VAR_in25;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_iffalse := VAR_in26;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_iftrue := VAR_in27;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_iffalse := VAR_in28;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_iftrue := VAR_in29;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_iftrue := VAR_in3;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_iffalse := VAR_in30;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_iftrue := VAR_in31;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_iffalse := VAR_in32;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_iftrue := VAR_in33;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iffalse := VAR_in34;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iftrue := VAR_in35;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_iffalse := VAR_in36;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_iftrue := VAR_in37;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_iffalse := VAR_in38;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_iftrue := VAR_in39;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_iffalse := VAR_in4;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_iffalse := VAR_in40;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_iftrue := VAR_in41;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_iffalse := VAR_in42;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_iftrue := VAR_in43;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_iffalse := VAR_in44;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_iftrue := VAR_in45;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_iffalse := VAR_in46;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_iftrue := VAR_in47;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_iffalse := VAR_in48;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_iftrue := VAR_in49;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_iftrue := VAR_in5;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iffalse := VAR_in50;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iftrue := VAR_in51;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_iffalse := VAR_in52;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_iftrue := VAR_in53;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_iffalse := VAR_in54;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_iftrue := VAR_in55;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_iffalse := VAR_in56;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_iftrue := VAR_in57;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_iffalse := VAR_in58;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_iftrue := VAR_in59;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_iffalse := VAR_in6;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iffalse := VAR_in60;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iftrue := VAR_in61;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_iffalse := VAR_in62;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_iftrue := VAR_in63;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_iffalse := VAR_in64;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_iftrue := VAR_in65;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_iffalse := VAR_in66;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_iftrue := VAR_in67;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_iffalse := VAR_in68;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_iftrue := VAR_in69;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_iftrue := VAR_in7;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_iffalse := VAR_in70;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_iftrue := VAR_in71;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_iffalse := VAR_in72;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_iftrue := VAR_in73;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_iffalse := VAR_in74;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_iftrue := VAR_in75;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iffalse := VAR_in76;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iftrue := VAR_in77;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_iffalse := VAR_in78;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_iftrue := VAR_in79;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_iffalse := VAR_in8;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_iffalse := VAR_in80;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_iftrue := VAR_in81;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_iffalse := VAR_in82;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_iftrue := VAR_in83;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_iffalse := VAR_in84;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_iftrue := VAR_in85;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iffalse := VAR_in86;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iftrue := VAR_in87;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_iffalse := VAR_in88;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_iftrue := VAR_in89;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_iftrue := VAR_in9;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_iffalse := VAR_in90;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_iftrue := VAR_in91;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_iffalse := VAR_in92;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_iftrue := VAR_in93;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_iffalse := VAR_in94;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_iftrue := VAR_in95;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iffalse := VAR_in96;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iftrue := VAR_in97;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_iffalse := VAR_in98;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_iftrue := VAR_in99;
     -- uint7_1_1[bit_math_h_l724_c10_6bba] LATENCY=0
     VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output := uint7_1_1(
     VAR_sel);

     -- uint7_4_4[bit_math_h_l1358_c10_7de3] LATENCY=0
     VAR_uint7_4_4_bit_math_h_l1358_c10_7de3_return_output := uint7_4_4(
     VAR_sel);

     -- uint7_3_3[bit_math_h_l1264_c10_0dc7] LATENCY=0
     VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output := uint7_3_3(
     VAR_sel);

     -- uint7_2_2[bit_math_h_l1082_c10_9337] LATENCY=0
     VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output := uint7_2_2(
     VAR_sel);

     -- uint7_0_0[bit_math_h_l14_c10_703d] LATENCY=0
     VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output := uint7_0_0(
     VAR_sel);

     -- uint7_5_5[bit_math_h_l1408_c10_6715] LATENCY=0
     VAR_uint7_5_5_bit_math_h_l1408_c10_6715_return_output := uint7_5_5(
     VAR_sel);

     -- uint7_6_6[bit_math_h_l1436_c10_2546] LATENCY=0
     VAR_uint7_6_6_bit_math_h_l1436_c10_2546_return_output := uint7_6_6(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_cond := VAR_uint7_0_0_bit_math_h_l14_c10_703d_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_cond := VAR_uint7_1_1_bit_math_h_l724_c10_6bba_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_9337_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_0dc7_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_7de3_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_7de3_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_7de3_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_7de3_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_6715_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_6715_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_cond := VAR_uint7_6_6_bit_math_h_l1436_c10_2546_return_output;
     -- layer0_node47_MUX[bit_math_h_l535_c3_18b2] LATENCY=0
     -- Inputs
     layer0_node47_MUX_bit_math_h_l535_c3_18b2_cond <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_cond;
     layer0_node47_MUX_bit_math_h_l535_c3_18b2_iftrue <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_iftrue;
     layer0_node47_MUX_bit_math_h_l535_c3_18b2_iffalse <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_iffalse;
     -- Outputs
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_return_output := layer0_node47_MUX_bit_math_h_l535_c3_18b2_return_output;

     -- layer0_node6_MUX[bit_math_h_l84_c3_494b] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_494b_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_494b_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_494b_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_return_output := layer0_node6_MUX_bit_math_h_l84_c3_494b_return_output;

     -- layer0_node27_MUX[bit_math_h_l315_c3_7789] LATENCY=0
     -- Inputs
     layer0_node27_MUX_bit_math_h_l315_c3_7789_cond <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_cond;
     layer0_node27_MUX_bit_math_h_l315_c3_7789_iftrue <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_iftrue;
     layer0_node27_MUX_bit_math_h_l315_c3_7789_iffalse <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_iffalse;
     -- Outputs
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_return_output := layer0_node27_MUX_bit_math_h_l315_c3_7789_return_output;

     -- layer0_node17_MUX[bit_math_h_l205_c3_4b2c] LATENCY=0
     -- Inputs
     layer0_node17_MUX_bit_math_h_l205_c3_4b2c_cond <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_cond;
     layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iftrue <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iftrue;
     layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iffalse <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_iffalse;
     -- Outputs
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_return_output := layer0_node17_MUX_bit_math_h_l205_c3_4b2c_return_output;

     -- layer0_node39_MUX[bit_math_h_l447_c3_7b35] LATENCY=0
     -- Inputs
     layer0_node39_MUX_bit_math_h_l447_c3_7b35_cond <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_cond;
     layer0_node39_MUX_bit_math_h_l447_c3_7b35_iftrue <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_iftrue;
     layer0_node39_MUX_bit_math_h_l447_c3_7b35_iffalse <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_iffalse;
     -- Outputs
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_return_output := layer0_node39_MUX_bit_math_h_l447_c3_7b35_return_output;

     -- layer0_node29_MUX[bit_math_h_l337_c3_9c87] LATENCY=0
     -- Inputs
     layer0_node29_MUX_bit_math_h_l337_c3_9c87_cond <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_cond;
     layer0_node29_MUX_bit_math_h_l337_c3_9c87_iftrue <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_iftrue;
     layer0_node29_MUX_bit_math_h_l337_c3_9c87_iffalse <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_iffalse;
     -- Outputs
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_return_output := layer0_node29_MUX_bit_math_h_l337_c3_9c87_return_output;

     -- layer0_node49_MUX[bit_math_h_l557_c3_68c1] LATENCY=0
     -- Inputs
     layer0_node49_MUX_bit_math_h_l557_c3_68c1_cond <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_cond;
     layer0_node49_MUX_bit_math_h_l557_c3_68c1_iftrue <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_iftrue;
     layer0_node49_MUX_bit_math_h_l557_c3_68c1_iffalse <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_iffalse;
     -- Outputs
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_return_output := layer0_node49_MUX_bit_math_h_l557_c3_68c1_return_output;

     -- layer0_node13_MUX[bit_math_h_l161_c3_c865] LATENCY=0
     -- Inputs
     layer0_node13_MUX_bit_math_h_l161_c3_c865_cond <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_cond;
     layer0_node13_MUX_bit_math_h_l161_c3_c865_iftrue <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_iftrue;
     layer0_node13_MUX_bit_math_h_l161_c3_c865_iffalse <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_iffalse;
     -- Outputs
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_return_output := layer0_node13_MUX_bit_math_h_l161_c3_c865_return_output;

     -- layer0_node61_MUX[bit_math_h_l689_c3_580e] LATENCY=0
     -- Inputs
     layer0_node61_MUX_bit_math_h_l689_c3_580e_cond <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_cond;
     layer0_node61_MUX_bit_math_h_l689_c3_580e_iftrue <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_iftrue;
     layer0_node61_MUX_bit_math_h_l689_c3_580e_iffalse <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_iffalse;
     -- Outputs
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_return_output := layer0_node61_MUX_bit_math_h_l689_c3_580e_return_output;

     -- layer0_node15_MUX[bit_math_h_l183_c3_6211] LATENCY=0
     -- Inputs
     layer0_node15_MUX_bit_math_h_l183_c3_6211_cond <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_cond;
     layer0_node15_MUX_bit_math_h_l183_c3_6211_iftrue <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_iftrue;
     layer0_node15_MUX_bit_math_h_l183_c3_6211_iffalse <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_iffalse;
     -- Outputs
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_return_output := layer0_node15_MUX_bit_math_h_l183_c3_6211_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_daab] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_daab_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_daab_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_daab_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_return_output := layer0_node7_MUX_bit_math_h_l95_c3_daab_return_output;

     -- layer0_node59_MUX[bit_math_h_l667_c3_b104] LATENCY=0
     -- Inputs
     layer0_node59_MUX_bit_math_h_l667_c3_b104_cond <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_cond;
     layer0_node59_MUX_bit_math_h_l667_c3_b104_iftrue <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_iftrue;
     layer0_node59_MUX_bit_math_h_l667_c3_b104_iffalse <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_iffalse;
     -- Outputs
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_return_output := layer0_node59_MUX_bit_math_h_l667_c3_b104_return_output;

     -- layer0_node60_MUX[bit_math_h_l678_c3_7571] LATENCY=0
     -- Inputs
     layer0_node60_MUX_bit_math_h_l678_c3_7571_cond <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_cond;
     layer0_node60_MUX_bit_math_h_l678_c3_7571_iftrue <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_iftrue;
     layer0_node60_MUX_bit_math_h_l678_c3_7571_iffalse <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_iffalse;
     -- Outputs
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_return_output := layer0_node60_MUX_bit_math_h_l678_c3_7571_return_output;

     -- layer0_node12_MUX[bit_math_h_l150_c3_af2c] LATENCY=0
     -- Inputs
     layer0_node12_MUX_bit_math_h_l150_c3_af2c_cond <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_cond;
     layer0_node12_MUX_bit_math_h_l150_c3_af2c_iftrue <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_iftrue;
     layer0_node12_MUX_bit_math_h_l150_c3_af2c_iffalse <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_iffalse;
     -- Outputs
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_return_output := layer0_node12_MUX_bit_math_h_l150_c3_af2c_return_output;

     -- layer0_node32_MUX[bit_math_h_l370_c3_4893] LATENCY=0
     -- Inputs
     layer0_node32_MUX_bit_math_h_l370_c3_4893_cond <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_cond;
     layer0_node32_MUX_bit_math_h_l370_c3_4893_iftrue <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_iftrue;
     layer0_node32_MUX_bit_math_h_l370_c3_4893_iffalse <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_iffalse;
     -- Outputs
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_return_output := layer0_node32_MUX_bit_math_h_l370_c3_4893_return_output;

     -- layer0_node10_MUX[bit_math_h_l128_c3_06d1] LATENCY=0
     -- Inputs
     layer0_node10_MUX_bit_math_h_l128_c3_06d1_cond <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_cond;
     layer0_node10_MUX_bit_math_h_l128_c3_06d1_iftrue <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_iftrue;
     layer0_node10_MUX_bit_math_h_l128_c3_06d1_iffalse <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_iffalse;
     -- Outputs
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_return_output := layer0_node10_MUX_bit_math_h_l128_c3_06d1_return_output;

     -- layer0_node1_MUX[bit_math_h_l29_c3_dc12] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_dc12_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_dc12_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_dc12_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_return_output := layer0_node1_MUX_bit_math_h_l29_c3_dc12_return_output;

     -- layer0_node18_MUX[bit_math_h_l216_c3_0b83] LATENCY=0
     -- Inputs
     layer0_node18_MUX_bit_math_h_l216_c3_0b83_cond <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_cond;
     layer0_node18_MUX_bit_math_h_l216_c3_0b83_iftrue <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_iftrue;
     layer0_node18_MUX_bit_math_h_l216_c3_0b83_iffalse <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_iffalse;
     -- Outputs
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_return_output := layer0_node18_MUX_bit_math_h_l216_c3_0b83_return_output;

     -- layer0_node36_MUX[bit_math_h_l414_c3_7348] LATENCY=0
     -- Inputs
     layer0_node36_MUX_bit_math_h_l414_c3_7348_cond <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_cond;
     layer0_node36_MUX_bit_math_h_l414_c3_7348_iftrue <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_iftrue;
     layer0_node36_MUX_bit_math_h_l414_c3_7348_iffalse <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_iffalse;
     -- Outputs
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_return_output := layer0_node36_MUX_bit_math_h_l414_c3_7348_return_output;

     -- layer0_node8_MUX[bit_math_h_l106_c3_d50d] LATENCY=0
     -- Inputs
     layer0_node8_MUX_bit_math_h_l106_c3_d50d_cond <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_cond;
     layer0_node8_MUX_bit_math_h_l106_c3_d50d_iftrue <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_iftrue;
     layer0_node8_MUX_bit_math_h_l106_c3_d50d_iffalse <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_iffalse;
     -- Outputs
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_return_output := layer0_node8_MUX_bit_math_h_l106_c3_d50d_return_output;

     -- layer0_node50_MUX[bit_math_h_l568_c3_8ec7] LATENCY=0
     -- Inputs
     layer0_node50_MUX_bit_math_h_l568_c3_8ec7_cond <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_cond;
     layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iftrue <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iftrue;
     layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iffalse <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_iffalse;
     -- Outputs
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_return_output := layer0_node50_MUX_bit_math_h_l568_c3_8ec7_return_output;

     -- layer0_node51_MUX[bit_math_h_l579_c3_5985] LATENCY=0
     -- Inputs
     layer0_node51_MUX_bit_math_h_l579_c3_5985_cond <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_cond;
     layer0_node51_MUX_bit_math_h_l579_c3_5985_iftrue <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_iftrue;
     layer0_node51_MUX_bit_math_h_l579_c3_5985_iffalse <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_iffalse;
     -- Outputs
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_return_output := layer0_node51_MUX_bit_math_h_l579_c3_5985_return_output;

     -- layer0_node44_MUX[bit_math_h_l502_c3_84a4] LATENCY=0
     -- Inputs
     layer0_node44_MUX_bit_math_h_l502_c3_84a4_cond <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_cond;
     layer0_node44_MUX_bit_math_h_l502_c3_84a4_iftrue <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_iftrue;
     layer0_node44_MUX_bit_math_h_l502_c3_84a4_iffalse <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_iffalse;
     -- Outputs
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_return_output := layer0_node44_MUX_bit_math_h_l502_c3_84a4_return_output;

     -- layer0_node38_MUX[bit_math_h_l436_c3_d3a0] LATENCY=0
     -- Inputs
     layer0_node38_MUX_bit_math_h_l436_c3_d3a0_cond <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_cond;
     layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iftrue <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iftrue;
     layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iffalse <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_iffalse;
     -- Outputs
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_return_output := layer0_node38_MUX_bit_math_h_l436_c3_d3a0_return_output;

     -- layer0_node34_MUX[bit_math_h_l392_c3_59bd] LATENCY=0
     -- Inputs
     layer0_node34_MUX_bit_math_h_l392_c3_59bd_cond <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_cond;
     layer0_node34_MUX_bit_math_h_l392_c3_59bd_iftrue <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_iftrue;
     layer0_node34_MUX_bit_math_h_l392_c3_59bd_iffalse <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_iffalse;
     -- Outputs
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_return_output := layer0_node34_MUX_bit_math_h_l392_c3_59bd_return_output;

     -- layer0_node9_MUX[bit_math_h_l117_c3_c9ee] LATENCY=0
     -- Inputs
     layer0_node9_MUX_bit_math_h_l117_c3_c9ee_cond <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_cond;
     layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iftrue <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iftrue;
     layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iffalse <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_iffalse;
     -- Outputs
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_return_output := layer0_node9_MUX_bit_math_h_l117_c3_c9ee_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_70c7] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_70c7_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_70c7_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_70c7_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_return_output := layer0_node0_MUX_bit_math_h_l18_c3_70c7_return_output;

     -- layer0_node25_MUX[bit_math_h_l293_c3_b4b9] LATENCY=0
     -- Inputs
     layer0_node25_MUX_bit_math_h_l293_c3_b4b9_cond <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_cond;
     layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iftrue <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iftrue;
     layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iffalse <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_iffalse;
     -- Outputs
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_return_output := layer0_node25_MUX_bit_math_h_l293_c3_b4b9_return_output;

     -- layer0_node28_MUX[bit_math_h_l326_c3_098d] LATENCY=0
     -- Inputs
     layer0_node28_MUX_bit_math_h_l326_c3_098d_cond <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_cond;
     layer0_node28_MUX_bit_math_h_l326_c3_098d_iftrue <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_iftrue;
     layer0_node28_MUX_bit_math_h_l326_c3_098d_iffalse <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_iffalse;
     -- Outputs
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_return_output := layer0_node28_MUX_bit_math_h_l326_c3_098d_return_output;

     -- layer0_node58_MUX[bit_math_h_l656_c3_b995] LATENCY=0
     -- Inputs
     layer0_node58_MUX_bit_math_h_l656_c3_b995_cond <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_cond;
     layer0_node58_MUX_bit_math_h_l656_c3_b995_iftrue <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_iftrue;
     layer0_node58_MUX_bit_math_h_l656_c3_b995_iffalse <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_iffalse;
     -- Outputs
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_return_output := layer0_node58_MUX_bit_math_h_l656_c3_b995_return_output;

     -- layer0_node46_MUX[bit_math_h_l524_c3_42cd] LATENCY=0
     -- Inputs
     layer0_node46_MUX_bit_math_h_l524_c3_42cd_cond <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_cond;
     layer0_node46_MUX_bit_math_h_l524_c3_42cd_iftrue <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_iftrue;
     layer0_node46_MUX_bit_math_h_l524_c3_42cd_iffalse <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_iffalse;
     -- Outputs
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_return_output := layer0_node46_MUX_bit_math_h_l524_c3_42cd_return_output;

     -- layer0_node21_MUX[bit_math_h_l249_c3_c173] LATENCY=0
     -- Inputs
     layer0_node21_MUX_bit_math_h_l249_c3_c173_cond <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_cond;
     layer0_node21_MUX_bit_math_h_l249_c3_c173_iftrue <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_iftrue;
     layer0_node21_MUX_bit_math_h_l249_c3_c173_iffalse <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_iffalse;
     -- Outputs
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_return_output := layer0_node21_MUX_bit_math_h_l249_c3_c173_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_3404] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_3404_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_3404_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_3404_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_return_output := layer0_node2_MUX_bit_math_h_l40_c3_3404_return_output;

     -- layer0_node26_MUX[bit_math_h_l304_c3_2bce] LATENCY=0
     -- Inputs
     layer0_node26_MUX_bit_math_h_l304_c3_2bce_cond <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_cond;
     layer0_node26_MUX_bit_math_h_l304_c3_2bce_iftrue <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_iftrue;
     layer0_node26_MUX_bit_math_h_l304_c3_2bce_iffalse <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_iffalse;
     -- Outputs
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_return_output := layer0_node26_MUX_bit_math_h_l304_c3_2bce_return_output;

     -- layer0_node45_MUX[bit_math_h_l513_c3_552e] LATENCY=0
     -- Inputs
     layer0_node45_MUX_bit_math_h_l513_c3_552e_cond <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_cond;
     layer0_node45_MUX_bit_math_h_l513_c3_552e_iftrue <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_iftrue;
     layer0_node45_MUX_bit_math_h_l513_c3_552e_iffalse <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_iffalse;
     -- Outputs
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_return_output := layer0_node45_MUX_bit_math_h_l513_c3_552e_return_output;

     -- layer0_node63_MUX[bit_math_h_l711_c3_17f2] LATENCY=0
     -- Inputs
     layer0_node63_MUX_bit_math_h_l711_c3_17f2_cond <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_cond;
     layer0_node63_MUX_bit_math_h_l711_c3_17f2_iftrue <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_iftrue;
     layer0_node63_MUX_bit_math_h_l711_c3_17f2_iffalse <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_iffalse;
     -- Outputs
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_return_output := layer0_node63_MUX_bit_math_h_l711_c3_17f2_return_output;

     -- layer0_node31_MUX[bit_math_h_l359_c3_5065] LATENCY=0
     -- Inputs
     layer0_node31_MUX_bit_math_h_l359_c3_5065_cond <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_cond;
     layer0_node31_MUX_bit_math_h_l359_c3_5065_iftrue <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_iftrue;
     layer0_node31_MUX_bit_math_h_l359_c3_5065_iffalse <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_iffalse;
     -- Outputs
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_return_output := layer0_node31_MUX_bit_math_h_l359_c3_5065_return_output;

     -- layer0_node19_MUX[bit_math_h_l227_c3_1e36] LATENCY=0
     -- Inputs
     layer0_node19_MUX_bit_math_h_l227_c3_1e36_cond <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_cond;
     layer0_node19_MUX_bit_math_h_l227_c3_1e36_iftrue <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_iftrue;
     layer0_node19_MUX_bit_math_h_l227_c3_1e36_iffalse <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_iffalse;
     -- Outputs
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_return_output := layer0_node19_MUX_bit_math_h_l227_c3_1e36_return_output;

     -- layer0_node48_MUX[bit_math_h_l546_c3_e9fe] LATENCY=0
     -- Inputs
     layer0_node48_MUX_bit_math_h_l546_c3_e9fe_cond <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_cond;
     layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iftrue <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iftrue;
     layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iffalse <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_iffalse;
     -- Outputs
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_return_output := layer0_node48_MUX_bit_math_h_l546_c3_e9fe_return_output;

     -- layer0_node43_MUX[bit_math_h_l491_c3_6ed7] LATENCY=0
     -- Inputs
     layer0_node43_MUX_bit_math_h_l491_c3_6ed7_cond <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_cond;
     layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iftrue <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iftrue;
     layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iffalse <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_iffalse;
     -- Outputs
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_return_output := layer0_node43_MUX_bit_math_h_l491_c3_6ed7_return_output;

     -- layer0_node30_MUX[bit_math_h_l348_c3_6b0d] LATENCY=0
     -- Inputs
     layer0_node30_MUX_bit_math_h_l348_c3_6b0d_cond <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_cond;
     layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iftrue <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iftrue;
     layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iffalse <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_iffalse;
     -- Outputs
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_return_output := layer0_node30_MUX_bit_math_h_l348_c3_6b0d_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_cc01] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_cc01_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_cc01_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_cc01_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_return_output := layer0_node3_MUX_bit_math_h_l51_c3_cc01_return_output;

     -- layer0_node52_MUX[bit_math_h_l590_c3_90c2] LATENCY=0
     -- Inputs
     layer0_node52_MUX_bit_math_h_l590_c3_90c2_cond <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_cond;
     layer0_node52_MUX_bit_math_h_l590_c3_90c2_iftrue <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_iftrue;
     layer0_node52_MUX_bit_math_h_l590_c3_90c2_iffalse <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_iffalse;
     -- Outputs
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_return_output := layer0_node52_MUX_bit_math_h_l590_c3_90c2_return_output;

     -- layer0_node41_MUX[bit_math_h_l469_c3_47d5] LATENCY=0
     -- Inputs
     layer0_node41_MUX_bit_math_h_l469_c3_47d5_cond <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_cond;
     layer0_node41_MUX_bit_math_h_l469_c3_47d5_iftrue <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_iftrue;
     layer0_node41_MUX_bit_math_h_l469_c3_47d5_iffalse <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_iffalse;
     -- Outputs
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_return_output := layer0_node41_MUX_bit_math_h_l469_c3_47d5_return_output;

     -- layer0_node22_MUX[bit_math_h_l260_c3_fce5] LATENCY=0
     -- Inputs
     layer0_node22_MUX_bit_math_h_l260_c3_fce5_cond <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_cond;
     layer0_node22_MUX_bit_math_h_l260_c3_fce5_iftrue <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_iftrue;
     layer0_node22_MUX_bit_math_h_l260_c3_fce5_iffalse <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_iffalse;
     -- Outputs
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_return_output := layer0_node22_MUX_bit_math_h_l260_c3_fce5_return_output;

     -- layer0_node53_MUX[bit_math_h_l601_c3_5a9e] LATENCY=0
     -- Inputs
     layer0_node53_MUX_bit_math_h_l601_c3_5a9e_cond <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_cond;
     layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iftrue <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iftrue;
     layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iffalse <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_iffalse;
     -- Outputs
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_return_output := layer0_node53_MUX_bit_math_h_l601_c3_5a9e_return_output;

     -- layer0_node57_MUX[bit_math_h_l645_c3_eeb0] LATENCY=0
     -- Inputs
     layer0_node57_MUX_bit_math_h_l645_c3_eeb0_cond <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_cond;
     layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iftrue <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iftrue;
     layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iffalse <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_iffalse;
     -- Outputs
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_return_output := layer0_node57_MUX_bit_math_h_l645_c3_eeb0_return_output;

     -- layer0_node23_MUX[bit_math_h_l271_c3_a82d] LATENCY=0
     -- Inputs
     layer0_node23_MUX_bit_math_h_l271_c3_a82d_cond <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_cond;
     layer0_node23_MUX_bit_math_h_l271_c3_a82d_iftrue <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_iftrue;
     layer0_node23_MUX_bit_math_h_l271_c3_a82d_iffalse <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_iffalse;
     -- Outputs
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_return_output := layer0_node23_MUX_bit_math_h_l271_c3_a82d_return_output;

     -- layer0_node56_MUX[bit_math_h_l634_c3_f6e3] LATENCY=0
     -- Inputs
     layer0_node56_MUX_bit_math_h_l634_c3_f6e3_cond <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_cond;
     layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iftrue <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iftrue;
     layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iffalse <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_iffalse;
     -- Outputs
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_return_output := layer0_node56_MUX_bit_math_h_l634_c3_f6e3_return_output;

     -- layer0_node16_MUX[bit_math_h_l194_c3_6e24] LATENCY=0
     -- Inputs
     layer0_node16_MUX_bit_math_h_l194_c3_6e24_cond <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_cond;
     layer0_node16_MUX_bit_math_h_l194_c3_6e24_iftrue <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_iftrue;
     layer0_node16_MUX_bit_math_h_l194_c3_6e24_iffalse <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_iffalse;
     -- Outputs
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_return_output := layer0_node16_MUX_bit_math_h_l194_c3_6e24_return_output;

     -- layer0_node5_MUX[bit_math_h_l73_c3_2acd] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_2acd_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_2acd_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_2acd_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_return_output := layer0_node5_MUX_bit_math_h_l73_c3_2acd_return_output;

     -- layer0_node37_MUX[bit_math_h_l425_c3_f929] LATENCY=0
     -- Inputs
     layer0_node37_MUX_bit_math_h_l425_c3_f929_cond <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_cond;
     layer0_node37_MUX_bit_math_h_l425_c3_f929_iftrue <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_iftrue;
     layer0_node37_MUX_bit_math_h_l425_c3_f929_iffalse <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_iffalse;
     -- Outputs
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_return_output := layer0_node37_MUX_bit_math_h_l425_c3_f929_return_output;

     -- layer0_node62_MUX[bit_math_h_l700_c3_9f5f] LATENCY=0
     -- Inputs
     layer0_node62_MUX_bit_math_h_l700_c3_9f5f_cond <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_cond;
     layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iftrue <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iftrue;
     layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iffalse <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_iffalse;
     -- Outputs
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_return_output := layer0_node62_MUX_bit_math_h_l700_c3_9f5f_return_output;

     -- layer0_node42_MUX[bit_math_h_l480_c3_50c3] LATENCY=0
     -- Inputs
     layer0_node42_MUX_bit_math_h_l480_c3_50c3_cond <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_cond;
     layer0_node42_MUX_bit_math_h_l480_c3_50c3_iftrue <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_iftrue;
     layer0_node42_MUX_bit_math_h_l480_c3_50c3_iffalse <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_iffalse;
     -- Outputs
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_return_output := layer0_node42_MUX_bit_math_h_l480_c3_50c3_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_7793] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_7793_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_7793_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_7793_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_return_output := layer0_node4_MUX_bit_math_h_l62_c3_7793_return_output;

     -- layer0_node11_MUX[bit_math_h_l139_c3_13dc] LATENCY=0
     -- Inputs
     layer0_node11_MUX_bit_math_h_l139_c3_13dc_cond <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_cond;
     layer0_node11_MUX_bit_math_h_l139_c3_13dc_iftrue <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_iftrue;
     layer0_node11_MUX_bit_math_h_l139_c3_13dc_iffalse <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_iffalse;
     -- Outputs
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_return_output := layer0_node11_MUX_bit_math_h_l139_c3_13dc_return_output;

     -- layer0_node20_MUX[bit_math_h_l238_c3_5458] LATENCY=0
     -- Inputs
     layer0_node20_MUX_bit_math_h_l238_c3_5458_cond <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_cond;
     layer0_node20_MUX_bit_math_h_l238_c3_5458_iftrue <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_iftrue;
     layer0_node20_MUX_bit_math_h_l238_c3_5458_iffalse <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_iffalse;
     -- Outputs
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_return_output := layer0_node20_MUX_bit_math_h_l238_c3_5458_return_output;

     -- layer0_node54_MUX[bit_math_h_l612_c3_235a] LATENCY=0
     -- Inputs
     layer0_node54_MUX_bit_math_h_l612_c3_235a_cond <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_cond;
     layer0_node54_MUX_bit_math_h_l612_c3_235a_iftrue <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_iftrue;
     layer0_node54_MUX_bit_math_h_l612_c3_235a_iffalse <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_iffalse;
     -- Outputs
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_return_output := layer0_node54_MUX_bit_math_h_l612_c3_235a_return_output;

     -- layer0_node24_MUX[bit_math_h_l282_c3_6611] LATENCY=0
     -- Inputs
     layer0_node24_MUX_bit_math_h_l282_c3_6611_cond <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_cond;
     layer0_node24_MUX_bit_math_h_l282_c3_6611_iftrue <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_iftrue;
     layer0_node24_MUX_bit_math_h_l282_c3_6611_iffalse <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_iffalse;
     -- Outputs
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_return_output := layer0_node24_MUX_bit_math_h_l282_c3_6611_return_output;

     -- layer0_node55_MUX[bit_math_h_l623_c3_1dea] LATENCY=0
     -- Inputs
     layer0_node55_MUX_bit_math_h_l623_c3_1dea_cond <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_cond;
     layer0_node55_MUX_bit_math_h_l623_c3_1dea_iftrue <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_iftrue;
     layer0_node55_MUX_bit_math_h_l623_c3_1dea_iffalse <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_iffalse;
     -- Outputs
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_return_output := layer0_node55_MUX_bit_math_h_l623_c3_1dea_return_output;

     -- layer0_node14_MUX[bit_math_h_l172_c3_1937] LATENCY=0
     -- Inputs
     layer0_node14_MUX_bit_math_h_l172_c3_1937_cond <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_cond;
     layer0_node14_MUX_bit_math_h_l172_c3_1937_iftrue <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_iftrue;
     layer0_node14_MUX_bit_math_h_l172_c3_1937_iffalse <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_iffalse;
     -- Outputs
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_return_output := layer0_node14_MUX_bit_math_h_l172_c3_1937_return_output;

     -- layer0_node33_MUX[bit_math_h_l381_c3_8132] LATENCY=0
     -- Inputs
     layer0_node33_MUX_bit_math_h_l381_c3_8132_cond <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_cond;
     layer0_node33_MUX_bit_math_h_l381_c3_8132_iftrue <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_iftrue;
     layer0_node33_MUX_bit_math_h_l381_c3_8132_iffalse <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_iffalse;
     -- Outputs
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_return_output := layer0_node33_MUX_bit_math_h_l381_c3_8132_return_output;

     -- layer0_node40_MUX[bit_math_h_l458_c3_426b] LATENCY=0
     -- Inputs
     layer0_node40_MUX_bit_math_h_l458_c3_426b_cond <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_cond;
     layer0_node40_MUX_bit_math_h_l458_c3_426b_iftrue <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_iftrue;
     layer0_node40_MUX_bit_math_h_l458_c3_426b_iffalse <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_iffalse;
     -- Outputs
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_return_output := layer0_node40_MUX_bit_math_h_l458_c3_426b_return_output;

     -- layer0_node35_MUX[bit_math_h_l403_c3_6326] LATENCY=0
     -- Inputs
     layer0_node35_MUX_bit_math_h_l403_c3_6326_cond <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_cond;
     layer0_node35_MUX_bit_math_h_l403_c3_6326_iftrue <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_iftrue;
     layer0_node35_MUX_bit_math_h_l403_c3_6326_iffalse <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_iffalse;
     -- Outputs
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_return_output := layer0_node35_MUX_bit_math_h_l403_c3_6326_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_70c7_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iffalse := VAR_layer0_node10_MUX_bit_math_h_l128_c3_06d1_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iftrue := VAR_layer0_node11_MUX_bit_math_h_l139_c3_13dc_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iffalse := VAR_layer0_node12_MUX_bit_math_h_l150_c3_af2c_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iftrue := VAR_layer0_node13_MUX_bit_math_h_l161_c3_c865_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_iffalse := VAR_layer0_node14_MUX_bit_math_h_l172_c3_1937_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_iftrue := VAR_layer0_node15_MUX_bit_math_h_l183_c3_6211_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_iffalse := VAR_layer0_node16_MUX_bit_math_h_l194_c3_6e24_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_iftrue := VAR_layer0_node17_MUX_bit_math_h_l205_c3_4b2c_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_iffalse := VAR_layer0_node18_MUX_bit_math_h_l216_c3_0b83_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_iftrue := VAR_layer0_node19_MUX_bit_math_h_l227_c3_1e36_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_dc12_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_iffalse := VAR_layer0_node20_MUX_bit_math_h_l238_c3_5458_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_iftrue := VAR_layer0_node21_MUX_bit_math_h_l249_c3_c173_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_iffalse := VAR_layer0_node22_MUX_bit_math_h_l260_c3_fce5_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_iftrue := VAR_layer0_node23_MUX_bit_math_h_l271_c3_a82d_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iffalse := VAR_layer0_node24_MUX_bit_math_h_l282_c3_6611_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iftrue := VAR_layer0_node25_MUX_bit_math_h_l293_c3_b4b9_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_iffalse := VAR_layer0_node26_MUX_bit_math_h_l304_c3_2bce_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_iftrue := VAR_layer0_node27_MUX_bit_math_h_l315_c3_7789_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iffalse := VAR_layer0_node28_MUX_bit_math_h_l326_c3_098d_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iftrue := VAR_layer0_node29_MUX_bit_math_h_l337_c3_9c87_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_3404_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_iffalse := VAR_layer0_node30_MUX_bit_math_h_l348_c3_6b0d_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_iftrue := VAR_layer0_node31_MUX_bit_math_h_l359_c3_5065_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iffalse := VAR_layer0_node32_MUX_bit_math_h_l370_c3_4893_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iftrue := VAR_layer0_node33_MUX_bit_math_h_l381_c3_8132_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iffalse := VAR_layer0_node34_MUX_bit_math_h_l392_c3_59bd_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iftrue := VAR_layer0_node35_MUX_bit_math_h_l403_c3_6326_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_iffalse := VAR_layer0_node36_MUX_bit_math_h_l414_c3_7348_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_iftrue := VAR_layer0_node37_MUX_bit_math_h_l425_c3_f929_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iffalse := VAR_layer0_node38_MUX_bit_math_h_l436_c3_d3a0_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iftrue := VAR_layer0_node39_MUX_bit_math_h_l447_c3_7b35_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_cc01_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_iffalse := VAR_layer0_node40_MUX_bit_math_h_l458_c3_426b_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_iftrue := VAR_layer0_node41_MUX_bit_math_h_l469_c3_47d5_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_iffalse := VAR_layer0_node42_MUX_bit_math_h_l480_c3_50c3_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_iftrue := VAR_layer0_node43_MUX_bit_math_h_l491_c3_6ed7_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iffalse := VAR_layer0_node44_MUX_bit_math_h_l502_c3_84a4_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iftrue := VAR_layer0_node45_MUX_bit_math_h_l513_c3_552e_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iffalse := VAR_layer0_node46_MUX_bit_math_h_l524_c3_42cd_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iftrue := VAR_layer0_node47_MUX_bit_math_h_l535_c3_18b2_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_iffalse := VAR_layer0_node48_MUX_bit_math_h_l546_c3_e9fe_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_iftrue := VAR_layer0_node49_MUX_bit_math_h_l557_c3_68c1_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_7793_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_iffalse := VAR_layer0_node50_MUX_bit_math_h_l568_c3_8ec7_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_iftrue := VAR_layer0_node51_MUX_bit_math_h_l579_c3_5985_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_iffalse := VAR_layer0_node52_MUX_bit_math_h_l590_c3_90c2_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_iftrue := VAR_layer0_node53_MUX_bit_math_h_l601_c3_5a9e_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iffalse := VAR_layer0_node54_MUX_bit_math_h_l612_c3_235a_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iftrue := VAR_layer0_node55_MUX_bit_math_h_l623_c3_1dea_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_iffalse := VAR_layer0_node56_MUX_bit_math_h_l634_c3_f6e3_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_iftrue := VAR_layer0_node57_MUX_bit_math_h_l645_c3_eeb0_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iffalse := VAR_layer0_node58_MUX_bit_math_h_l656_c3_b995_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iftrue := VAR_layer0_node59_MUX_bit_math_h_l667_c3_b104_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_2acd_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iffalse := VAR_layer0_node60_MUX_bit_math_h_l678_c3_7571_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iftrue := VAR_layer0_node61_MUX_bit_math_h_l689_c3_580e_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iffalse := VAR_layer0_node62_MUX_bit_math_h_l700_c3_9f5f_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iftrue := VAR_layer0_node63_MUX_bit_math_h_l711_c3_17f2_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_494b_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_daab_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_iffalse := VAR_layer0_node8_MUX_bit_math_h_l106_c3_d50d_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_iftrue := VAR_layer0_node9_MUX_bit_math_h_l117_c3_c9ee_return_output;
     -- layer1_node28_MUX[bit_math_h_l1036_c3_d560] LATENCY=0
     -- Inputs
     layer1_node28_MUX_bit_math_h_l1036_c3_d560_cond <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_cond;
     layer1_node28_MUX_bit_math_h_l1036_c3_d560_iftrue <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_iftrue;
     layer1_node28_MUX_bit_math_h_l1036_c3_d560_iffalse <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_iffalse;
     -- Outputs
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_return_output := layer1_node28_MUX_bit_math_h_l1036_c3_d560_return_output;

     -- layer1_node11_MUX[bit_math_h_l849_c3_c418] LATENCY=0
     -- Inputs
     layer1_node11_MUX_bit_math_h_l849_c3_c418_cond <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_cond;
     layer1_node11_MUX_bit_math_h_l849_c3_c418_iftrue <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_iftrue;
     layer1_node11_MUX_bit_math_h_l849_c3_c418_iffalse <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_iffalse;
     -- Outputs
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_return_output := layer1_node11_MUX_bit_math_h_l849_c3_c418_return_output;

     -- layer1_node6_MUX[bit_math_h_l794_c3_f4dd] LATENCY=0
     -- Inputs
     layer1_node6_MUX_bit_math_h_l794_c3_f4dd_cond <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_cond;
     layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iftrue <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iftrue;
     layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iffalse <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_iffalse;
     -- Outputs
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_return_output := layer1_node6_MUX_bit_math_h_l794_c3_f4dd_return_output;

     -- layer1_node29_MUX[bit_math_h_l1047_c3_9f00] LATENCY=0
     -- Inputs
     layer1_node29_MUX_bit_math_h_l1047_c3_9f00_cond <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_cond;
     layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iftrue <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iftrue;
     layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iffalse <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_iffalse;
     -- Outputs
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_return_output := layer1_node29_MUX_bit_math_h_l1047_c3_9f00_return_output;

     -- layer1_node25_MUX[bit_math_h_l1003_c3_371a] LATENCY=0
     -- Inputs
     layer1_node25_MUX_bit_math_h_l1003_c3_371a_cond <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_cond;
     layer1_node25_MUX_bit_math_h_l1003_c3_371a_iftrue <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_iftrue;
     layer1_node25_MUX_bit_math_h_l1003_c3_371a_iffalse <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_iffalse;
     -- Outputs
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_return_output := layer1_node25_MUX_bit_math_h_l1003_c3_371a_return_output;

     -- layer1_node7_MUX[bit_math_h_l805_c3_e535] LATENCY=0
     -- Inputs
     layer1_node7_MUX_bit_math_h_l805_c3_e535_cond <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_cond;
     layer1_node7_MUX_bit_math_h_l805_c3_e535_iftrue <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_iftrue;
     layer1_node7_MUX_bit_math_h_l805_c3_e535_iffalse <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_iffalse;
     -- Outputs
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_return_output := layer1_node7_MUX_bit_math_h_l805_c3_e535_return_output;

     -- layer1_node18_MUX[bit_math_h_l926_c3_15bb] LATENCY=0
     -- Inputs
     layer1_node18_MUX_bit_math_h_l926_c3_15bb_cond <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_cond;
     layer1_node18_MUX_bit_math_h_l926_c3_15bb_iftrue <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_iftrue;
     layer1_node18_MUX_bit_math_h_l926_c3_15bb_iffalse <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_iffalse;
     -- Outputs
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_return_output := layer1_node18_MUX_bit_math_h_l926_c3_15bb_return_output;

     -- layer1_node19_MUX[bit_math_h_l937_c3_3ad6] LATENCY=0
     -- Inputs
     layer1_node19_MUX_bit_math_h_l937_c3_3ad6_cond <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_cond;
     layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iftrue <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iftrue;
     layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iffalse <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_iffalse;
     -- Outputs
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_return_output := layer1_node19_MUX_bit_math_h_l937_c3_3ad6_return_output;

     -- layer1_node14_MUX[bit_math_h_l882_c3_5e4a] LATENCY=0
     -- Inputs
     layer1_node14_MUX_bit_math_h_l882_c3_5e4a_cond <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_cond;
     layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iftrue <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iftrue;
     layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iffalse <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_iffalse;
     -- Outputs
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_return_output := layer1_node14_MUX_bit_math_h_l882_c3_5e4a_return_output;

     -- layer1_node26_MUX[bit_math_h_l1014_c3_b858] LATENCY=0
     -- Inputs
     layer1_node26_MUX_bit_math_h_l1014_c3_b858_cond <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_cond;
     layer1_node26_MUX_bit_math_h_l1014_c3_b858_iftrue <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_iftrue;
     layer1_node26_MUX_bit_math_h_l1014_c3_b858_iffalse <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_iffalse;
     -- Outputs
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_return_output := layer1_node26_MUX_bit_math_h_l1014_c3_b858_return_output;

     -- layer1_node1_MUX[bit_math_h_l739_c3_57f6] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l739_c3_57f6_cond <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_cond;
     layer1_node1_MUX_bit_math_h_l739_c3_57f6_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_iftrue;
     layer1_node1_MUX_bit_math_h_l739_c3_57f6_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_return_output := layer1_node1_MUX_bit_math_h_l739_c3_57f6_return_output;

     -- layer1_node8_MUX[bit_math_h_l816_c3_e51d] LATENCY=0
     -- Inputs
     layer1_node8_MUX_bit_math_h_l816_c3_e51d_cond <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_cond;
     layer1_node8_MUX_bit_math_h_l816_c3_e51d_iftrue <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_iftrue;
     layer1_node8_MUX_bit_math_h_l816_c3_e51d_iffalse <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_iffalse;
     -- Outputs
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_return_output := layer1_node8_MUX_bit_math_h_l816_c3_e51d_return_output;

     -- layer1_node15_MUX[bit_math_h_l893_c3_faee] LATENCY=0
     -- Inputs
     layer1_node15_MUX_bit_math_h_l893_c3_faee_cond <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_cond;
     layer1_node15_MUX_bit_math_h_l893_c3_faee_iftrue <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_iftrue;
     layer1_node15_MUX_bit_math_h_l893_c3_faee_iffalse <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_iffalse;
     -- Outputs
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_return_output := layer1_node15_MUX_bit_math_h_l893_c3_faee_return_output;

     -- layer1_node17_MUX[bit_math_h_l915_c3_bbc7] LATENCY=0
     -- Inputs
     layer1_node17_MUX_bit_math_h_l915_c3_bbc7_cond <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_cond;
     layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iftrue <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iftrue;
     layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iffalse <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_iffalse;
     -- Outputs
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_return_output := layer1_node17_MUX_bit_math_h_l915_c3_bbc7_return_output;

     -- layer1_node5_MUX[bit_math_h_l783_c3_f8bc] LATENCY=0
     -- Inputs
     layer1_node5_MUX_bit_math_h_l783_c3_f8bc_cond <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_cond;
     layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iftrue <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iftrue;
     layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iffalse <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_iffalse;
     -- Outputs
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_return_output := layer1_node5_MUX_bit_math_h_l783_c3_f8bc_return_output;

     -- layer1_node27_MUX[bit_math_h_l1025_c3_d07c] LATENCY=0
     -- Inputs
     layer1_node27_MUX_bit_math_h_l1025_c3_d07c_cond <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_cond;
     layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iftrue <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iftrue;
     layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iffalse <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_iffalse;
     -- Outputs
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_return_output := layer1_node27_MUX_bit_math_h_l1025_c3_d07c_return_output;

     -- layer1_node23_MUX[bit_math_h_l981_c3_c1f3] LATENCY=0
     -- Inputs
     layer1_node23_MUX_bit_math_h_l981_c3_c1f3_cond <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_cond;
     layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iftrue <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iftrue;
     layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iffalse <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_iffalse;
     -- Outputs
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_return_output := layer1_node23_MUX_bit_math_h_l981_c3_c1f3_return_output;

     -- layer1_node4_MUX[bit_math_h_l772_c3_857f] LATENCY=0
     -- Inputs
     layer1_node4_MUX_bit_math_h_l772_c3_857f_cond <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_cond;
     layer1_node4_MUX_bit_math_h_l772_c3_857f_iftrue <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_iftrue;
     layer1_node4_MUX_bit_math_h_l772_c3_857f_iffalse <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_iffalse;
     -- Outputs
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_return_output := layer1_node4_MUX_bit_math_h_l772_c3_857f_return_output;

     -- layer1_node16_MUX[bit_math_h_l904_c3_1e1f] LATENCY=0
     -- Inputs
     layer1_node16_MUX_bit_math_h_l904_c3_1e1f_cond <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_cond;
     layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iftrue <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iftrue;
     layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iffalse <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_iffalse;
     -- Outputs
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_return_output := layer1_node16_MUX_bit_math_h_l904_c3_1e1f_return_output;

     -- layer1_node12_MUX[bit_math_h_l860_c3_3ea5] LATENCY=0
     -- Inputs
     layer1_node12_MUX_bit_math_h_l860_c3_3ea5_cond <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_cond;
     layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iftrue <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iftrue;
     layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iffalse <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_iffalse;
     -- Outputs
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_return_output := layer1_node12_MUX_bit_math_h_l860_c3_3ea5_return_output;

     -- layer1_node2_MUX[bit_math_h_l750_c3_b86b] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l750_c3_b86b_cond <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_cond;
     layer1_node2_MUX_bit_math_h_l750_c3_b86b_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_iftrue;
     layer1_node2_MUX_bit_math_h_l750_c3_b86b_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_return_output := layer1_node2_MUX_bit_math_h_l750_c3_b86b_return_output;

     -- layer1_node24_MUX[bit_math_h_l992_c3_1884] LATENCY=0
     -- Inputs
     layer1_node24_MUX_bit_math_h_l992_c3_1884_cond <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_cond;
     layer1_node24_MUX_bit_math_h_l992_c3_1884_iftrue <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_iftrue;
     layer1_node24_MUX_bit_math_h_l992_c3_1884_iffalse <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_iffalse;
     -- Outputs
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_return_output := layer1_node24_MUX_bit_math_h_l992_c3_1884_return_output;

     -- layer1_node9_MUX[bit_math_h_l827_c3_4f17] LATENCY=0
     -- Inputs
     layer1_node9_MUX_bit_math_h_l827_c3_4f17_cond <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_cond;
     layer1_node9_MUX_bit_math_h_l827_c3_4f17_iftrue <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_iftrue;
     layer1_node9_MUX_bit_math_h_l827_c3_4f17_iffalse <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_iffalse;
     -- Outputs
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_return_output := layer1_node9_MUX_bit_math_h_l827_c3_4f17_return_output;

     -- layer1_node21_MUX[bit_math_h_l959_c3_0003] LATENCY=0
     -- Inputs
     layer1_node21_MUX_bit_math_h_l959_c3_0003_cond <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_cond;
     layer1_node21_MUX_bit_math_h_l959_c3_0003_iftrue <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_iftrue;
     layer1_node21_MUX_bit_math_h_l959_c3_0003_iffalse <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_iffalse;
     -- Outputs
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_return_output := layer1_node21_MUX_bit_math_h_l959_c3_0003_return_output;

     -- layer1_node30_MUX[bit_math_h_l1058_c3_e6cc] LATENCY=0
     -- Inputs
     layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_cond <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_cond;
     layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iftrue <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iftrue;
     layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iffalse <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_iffalse;
     -- Outputs
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_return_output := layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_return_output;

     -- layer1_node3_MUX[bit_math_h_l761_c3_2586] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l761_c3_2586_cond <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_cond;
     layer1_node3_MUX_bit_math_h_l761_c3_2586_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_iftrue;
     layer1_node3_MUX_bit_math_h_l761_c3_2586_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_return_output := layer1_node3_MUX_bit_math_h_l761_c3_2586_return_output;

     -- layer1_node10_MUX[bit_math_h_l838_c3_8caa] LATENCY=0
     -- Inputs
     layer1_node10_MUX_bit_math_h_l838_c3_8caa_cond <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_cond;
     layer1_node10_MUX_bit_math_h_l838_c3_8caa_iftrue <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_iftrue;
     layer1_node10_MUX_bit_math_h_l838_c3_8caa_iffalse <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_iffalse;
     -- Outputs
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_return_output := layer1_node10_MUX_bit_math_h_l838_c3_8caa_return_output;

     -- layer1_node13_MUX[bit_math_h_l871_c3_66e4] LATENCY=0
     -- Inputs
     layer1_node13_MUX_bit_math_h_l871_c3_66e4_cond <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_cond;
     layer1_node13_MUX_bit_math_h_l871_c3_66e4_iftrue <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_iftrue;
     layer1_node13_MUX_bit_math_h_l871_c3_66e4_iffalse <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_iffalse;
     -- Outputs
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_return_output := layer1_node13_MUX_bit_math_h_l871_c3_66e4_return_output;

     -- layer1_node0_MUX[bit_math_h_l728_c3_23e3] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l728_c3_23e3_cond <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_cond;
     layer1_node0_MUX_bit_math_h_l728_c3_23e3_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_iftrue;
     layer1_node0_MUX_bit_math_h_l728_c3_23e3_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_return_output := layer1_node0_MUX_bit_math_h_l728_c3_23e3_return_output;

     -- layer1_node22_MUX[bit_math_h_l970_c3_fb2c] LATENCY=0
     -- Inputs
     layer1_node22_MUX_bit_math_h_l970_c3_fb2c_cond <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_cond;
     layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iftrue <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iftrue;
     layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iffalse <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_iffalse;
     -- Outputs
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_return_output := layer1_node22_MUX_bit_math_h_l970_c3_fb2c_return_output;

     -- layer1_node31_MUX[bit_math_h_l1069_c3_b1c7] LATENCY=0
     -- Inputs
     layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_cond <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_cond;
     layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iftrue <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iftrue;
     layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iffalse <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_iffalse;
     -- Outputs
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_return_output := layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_return_output;

     -- layer1_node20_MUX[bit_math_h_l948_c3_d497] LATENCY=0
     -- Inputs
     layer1_node20_MUX_bit_math_h_l948_c3_d497_cond <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_cond;
     layer1_node20_MUX_bit_math_h_l948_c3_d497_iftrue <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_iftrue;
     layer1_node20_MUX_bit_math_h_l948_c3_d497_iffalse <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_iffalse;
     -- Outputs
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_return_output := layer1_node20_MUX_bit_math_h_l948_c3_d497_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iffalse := VAR_layer1_node0_MUX_bit_math_h_l728_c3_23e3_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_iffalse := VAR_layer1_node10_MUX_bit_math_h_l838_c3_8caa_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_iftrue := VAR_layer1_node11_MUX_bit_math_h_l849_c3_c418_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iffalse := VAR_layer1_node12_MUX_bit_math_h_l860_c3_3ea5_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iftrue := VAR_layer1_node13_MUX_bit_math_h_l871_c3_66e4_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iffalse := VAR_layer1_node14_MUX_bit_math_h_l882_c3_5e4a_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iftrue := VAR_layer1_node15_MUX_bit_math_h_l893_c3_faee_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iffalse := VAR_layer1_node16_MUX_bit_math_h_l904_c3_1e1f_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iftrue := VAR_layer1_node17_MUX_bit_math_h_l915_c3_bbc7_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_iffalse := VAR_layer1_node18_MUX_bit_math_h_l926_c3_15bb_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_iftrue := VAR_layer1_node19_MUX_bit_math_h_l937_c3_3ad6_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iftrue := VAR_layer1_node1_MUX_bit_math_h_l739_c3_57f6_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_iffalse := VAR_layer1_node20_MUX_bit_math_h_l948_c3_d497_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_iftrue := VAR_layer1_node21_MUX_bit_math_h_l959_c3_0003_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iffalse := VAR_layer1_node22_MUX_bit_math_h_l970_c3_fb2c_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iftrue := VAR_layer1_node23_MUX_bit_math_h_l981_c3_c1f3_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iffalse := VAR_layer1_node24_MUX_bit_math_h_l992_c3_1884_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iftrue := VAR_layer1_node25_MUX_bit_math_h_l1003_c3_371a_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iffalse := VAR_layer1_node26_MUX_bit_math_h_l1014_c3_b858_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iftrue := VAR_layer1_node27_MUX_bit_math_h_l1025_c3_d07c_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iffalse := VAR_layer1_node28_MUX_bit_math_h_l1036_c3_d560_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iftrue := VAR_layer1_node29_MUX_bit_math_h_l1047_c3_9f00_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_iffalse := VAR_layer1_node2_MUX_bit_math_h_l750_c3_b86b_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iffalse := VAR_layer1_node30_MUX_bit_math_h_l1058_c3_e6cc_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iftrue := VAR_layer1_node31_MUX_bit_math_h_l1069_c3_b1c7_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_iftrue := VAR_layer1_node3_MUX_bit_math_h_l761_c3_2586_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iffalse := VAR_layer1_node4_MUX_bit_math_h_l772_c3_857f_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iftrue := VAR_layer1_node5_MUX_bit_math_h_l783_c3_f8bc_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_iffalse := VAR_layer1_node6_MUX_bit_math_h_l794_c3_f4dd_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_iftrue := VAR_layer1_node7_MUX_bit_math_h_l805_c3_e535_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_iffalse := VAR_layer1_node8_MUX_bit_math_h_l816_c3_e51d_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_iftrue := VAR_layer1_node9_MUX_bit_math_h_l827_c3_4f17_return_output;
     -- layer2_node1_MUX[bit_math_h_l1097_c3_7335] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l1097_c3_7335_cond <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_cond;
     layer2_node1_MUX_bit_math_h_l1097_c3_7335_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_iftrue;
     layer2_node1_MUX_bit_math_h_l1097_c3_7335_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_return_output := layer2_node1_MUX_bit_math_h_l1097_c3_7335_return_output;

     -- layer2_node13_MUX[bit_math_h_l1229_c3_bcb9] LATENCY=0
     -- Inputs
     layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_cond <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_cond;
     layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iftrue <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iftrue;
     layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iffalse <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_iffalse;
     -- Outputs
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_return_output := layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_return_output;

     -- layer2_node15_MUX[bit_math_h_l1251_c3_1e63] LATENCY=0
     -- Inputs
     layer2_node15_MUX_bit_math_h_l1251_c3_1e63_cond <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_cond;
     layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iftrue <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iftrue;
     layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iffalse <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_iffalse;
     -- Outputs
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_return_output := layer2_node15_MUX_bit_math_h_l1251_c3_1e63_return_output;

     -- layer2_node10_MUX[bit_math_h_l1196_c3_c187] LATENCY=0
     -- Inputs
     layer2_node10_MUX_bit_math_h_l1196_c3_c187_cond <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_cond;
     layer2_node10_MUX_bit_math_h_l1196_c3_c187_iftrue <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_iftrue;
     layer2_node10_MUX_bit_math_h_l1196_c3_c187_iffalse <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_iffalse;
     -- Outputs
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_return_output := layer2_node10_MUX_bit_math_h_l1196_c3_c187_return_output;

     -- layer2_node0_MUX[bit_math_h_l1086_c3_f3d3] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_cond <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_cond;
     layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iftrue;
     layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_return_output := layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_return_output;

     -- layer2_node6_MUX[bit_math_h_l1152_c3_be4a] LATENCY=0
     -- Inputs
     layer2_node6_MUX_bit_math_h_l1152_c3_be4a_cond <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_cond;
     layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iftrue <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iftrue;
     layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iffalse <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_iffalse;
     -- Outputs
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_return_output := layer2_node6_MUX_bit_math_h_l1152_c3_be4a_return_output;

     -- layer2_node11_MUX[bit_math_h_l1207_c3_bafc] LATENCY=0
     -- Inputs
     layer2_node11_MUX_bit_math_h_l1207_c3_bafc_cond <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_cond;
     layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iftrue <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iftrue;
     layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iffalse <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_iffalse;
     -- Outputs
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_return_output := layer2_node11_MUX_bit_math_h_l1207_c3_bafc_return_output;

     -- layer2_node9_MUX[bit_math_h_l1185_c3_e581] LATENCY=0
     -- Inputs
     layer2_node9_MUX_bit_math_h_l1185_c3_e581_cond <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_cond;
     layer2_node9_MUX_bit_math_h_l1185_c3_e581_iftrue <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_iftrue;
     layer2_node9_MUX_bit_math_h_l1185_c3_e581_iffalse <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_iffalse;
     -- Outputs
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_return_output := layer2_node9_MUX_bit_math_h_l1185_c3_e581_return_output;

     -- layer2_node14_MUX[bit_math_h_l1240_c3_7be3] LATENCY=0
     -- Inputs
     layer2_node14_MUX_bit_math_h_l1240_c3_7be3_cond <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_cond;
     layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iftrue <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iftrue;
     layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iffalse <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_iffalse;
     -- Outputs
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_return_output := layer2_node14_MUX_bit_math_h_l1240_c3_7be3_return_output;

     -- layer2_node4_MUX[bit_math_h_l1130_c3_0608] LATENCY=0
     -- Inputs
     layer2_node4_MUX_bit_math_h_l1130_c3_0608_cond <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_cond;
     layer2_node4_MUX_bit_math_h_l1130_c3_0608_iftrue <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_iftrue;
     layer2_node4_MUX_bit_math_h_l1130_c3_0608_iffalse <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_iffalse;
     -- Outputs
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_return_output := layer2_node4_MUX_bit_math_h_l1130_c3_0608_return_output;

     -- layer2_node7_MUX[bit_math_h_l1163_c3_4bab] LATENCY=0
     -- Inputs
     layer2_node7_MUX_bit_math_h_l1163_c3_4bab_cond <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_cond;
     layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iftrue <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iftrue;
     layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iffalse <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_iffalse;
     -- Outputs
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_return_output := layer2_node7_MUX_bit_math_h_l1163_c3_4bab_return_output;

     -- layer2_node8_MUX[bit_math_h_l1174_c3_24ff] LATENCY=0
     -- Inputs
     layer2_node8_MUX_bit_math_h_l1174_c3_24ff_cond <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_cond;
     layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iftrue <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iftrue;
     layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iffalse <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_iffalse;
     -- Outputs
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_return_output := layer2_node8_MUX_bit_math_h_l1174_c3_24ff_return_output;

     -- layer2_node12_MUX[bit_math_h_l1218_c3_c26f] LATENCY=0
     -- Inputs
     layer2_node12_MUX_bit_math_h_l1218_c3_c26f_cond <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_cond;
     layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iftrue <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iftrue;
     layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iffalse <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_iffalse;
     -- Outputs
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_return_output := layer2_node12_MUX_bit_math_h_l1218_c3_c26f_return_output;

     -- layer2_node2_MUX[bit_math_h_l1108_c3_bb5a] LATENCY=0
     -- Inputs
     layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_cond <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_cond;
     layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iftrue <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iftrue;
     layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iffalse <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_iffalse;
     -- Outputs
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_return_output := layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_return_output;

     -- layer2_node3_MUX[bit_math_h_l1119_c3_95be] LATENCY=0
     -- Inputs
     layer2_node3_MUX_bit_math_h_l1119_c3_95be_cond <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_cond;
     layer2_node3_MUX_bit_math_h_l1119_c3_95be_iftrue <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_iftrue;
     layer2_node3_MUX_bit_math_h_l1119_c3_95be_iffalse <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_iffalse;
     -- Outputs
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_return_output := layer2_node3_MUX_bit_math_h_l1119_c3_95be_return_output;

     -- layer2_node5_MUX[bit_math_h_l1141_c3_a965] LATENCY=0
     -- Inputs
     layer2_node5_MUX_bit_math_h_l1141_c3_a965_cond <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_cond;
     layer2_node5_MUX_bit_math_h_l1141_c3_a965_iftrue <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_iftrue;
     layer2_node5_MUX_bit_math_h_l1141_c3_a965_iffalse <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_iffalse;
     -- Outputs
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_return_output := layer2_node5_MUX_bit_math_h_l1141_c3_a965_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_iffalse := VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f3d3_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iffalse := VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c187_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iftrue := VAR_layer2_node11_MUX_bit_math_h_l1207_c3_bafc_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_iffalse := VAR_layer2_node12_MUX_bit_math_h_l1218_c3_c26f_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_iftrue := VAR_layer2_node13_MUX_bit_math_h_l1229_c3_bcb9_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iffalse := VAR_layer2_node14_MUX_bit_math_h_l1240_c3_7be3_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iftrue := VAR_layer2_node15_MUX_bit_math_h_l1251_c3_1e63_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_iftrue := VAR_layer2_node1_MUX_bit_math_h_l1097_c3_7335_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_iffalse := VAR_layer2_node2_MUX_bit_math_h_l1108_c3_bb5a_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_iftrue := VAR_layer2_node3_MUX_bit_math_h_l1119_c3_95be_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iffalse := VAR_layer2_node4_MUX_bit_math_h_l1130_c3_0608_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iftrue := VAR_layer2_node5_MUX_bit_math_h_l1141_c3_a965_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iffalse := VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be4a_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iftrue := VAR_layer2_node7_MUX_bit_math_h_l1163_c3_4bab_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_iffalse := VAR_layer2_node8_MUX_bit_math_h_l1174_c3_24ff_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_iftrue := VAR_layer2_node9_MUX_bit_math_h_l1185_c3_e581_return_output;
     -- layer3_node0_MUX[bit_math_h_l1268_c3_e356] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l1268_c3_e356_cond <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_cond;
     layer3_node0_MUX_bit_math_h_l1268_c3_e356_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_iftrue;
     layer3_node0_MUX_bit_math_h_l1268_c3_e356_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_return_output := layer3_node0_MUX_bit_math_h_l1268_c3_e356_return_output;

     -- layer3_node7_MUX[bit_math_h_l1345_c3_3cb2] LATENCY=0
     -- Inputs
     layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_cond <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_cond;
     layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iftrue <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iftrue;
     layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iffalse <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_iffalse;
     -- Outputs
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_return_output := layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_return_output;

     -- layer3_node1_MUX[bit_math_h_l1279_c3_3873] LATENCY=0
     -- Inputs
     layer3_node1_MUX_bit_math_h_l1279_c3_3873_cond <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_cond;
     layer3_node1_MUX_bit_math_h_l1279_c3_3873_iftrue <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_iftrue;
     layer3_node1_MUX_bit_math_h_l1279_c3_3873_iffalse <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_iffalse;
     -- Outputs
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_return_output := layer3_node1_MUX_bit_math_h_l1279_c3_3873_return_output;

     -- layer3_node2_MUX[bit_math_h_l1290_c3_4ec7] LATENCY=0
     -- Inputs
     layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_cond <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_cond;
     layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iftrue <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iftrue;
     layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iffalse <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_iffalse;
     -- Outputs
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_return_output := layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_return_output;

     -- layer3_node6_MUX[bit_math_h_l1334_c3_5def] LATENCY=0
     -- Inputs
     layer3_node6_MUX_bit_math_h_l1334_c3_5def_cond <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_cond;
     layer3_node6_MUX_bit_math_h_l1334_c3_5def_iftrue <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_iftrue;
     layer3_node6_MUX_bit_math_h_l1334_c3_5def_iffalse <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_iffalse;
     -- Outputs
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_return_output := layer3_node6_MUX_bit_math_h_l1334_c3_5def_return_output;

     -- layer3_node5_MUX[bit_math_h_l1323_c3_e63b] LATENCY=0
     -- Inputs
     layer3_node5_MUX_bit_math_h_l1323_c3_e63b_cond <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_cond;
     layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iftrue <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iftrue;
     layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iffalse <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_iffalse;
     -- Outputs
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_return_output := layer3_node5_MUX_bit_math_h_l1323_c3_e63b_return_output;

     -- layer3_node3_MUX[bit_math_h_l1301_c3_29f9] LATENCY=0
     -- Inputs
     layer3_node3_MUX_bit_math_h_l1301_c3_29f9_cond <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_cond;
     layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iftrue <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iftrue;
     layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iffalse <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_iffalse;
     -- Outputs
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_return_output := layer3_node3_MUX_bit_math_h_l1301_c3_29f9_return_output;

     -- layer3_node4_MUX[bit_math_h_l1312_c3_b484] LATENCY=0
     -- Inputs
     layer3_node4_MUX_bit_math_h_l1312_c3_b484_cond <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_cond;
     layer3_node4_MUX_bit_math_h_l1312_c3_b484_iftrue <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_iftrue;
     layer3_node4_MUX_bit_math_h_l1312_c3_b484_iffalse <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_iffalse;
     -- Outputs
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_return_output := layer3_node4_MUX_bit_math_h_l1312_c3_b484_return_output;

     -- Submodule level 5
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iffalse := VAR_layer3_node0_MUX_bit_math_h_l1268_c3_e356_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iftrue := VAR_layer3_node1_MUX_bit_math_h_l1279_c3_3873_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_iffalse := VAR_layer3_node2_MUX_bit_math_h_l1290_c3_4ec7_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_iftrue := VAR_layer3_node3_MUX_bit_math_h_l1301_c3_29f9_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_iffalse := VAR_layer3_node4_MUX_bit_math_h_l1312_c3_b484_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_iftrue := VAR_layer3_node5_MUX_bit_math_h_l1323_c3_e63b_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iffalse := VAR_layer3_node6_MUX_bit_math_h_l1334_c3_5def_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iftrue := VAR_layer3_node7_MUX_bit_math_h_l1345_c3_3cb2_return_output;
     -- layer4_node3_MUX[bit_math_h_l1395_c3_68f4] LATENCY=0
     -- Inputs
     layer4_node3_MUX_bit_math_h_l1395_c3_68f4_cond <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_cond;
     layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iftrue <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iftrue;
     layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iffalse <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_iffalse;
     -- Outputs
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_return_output := layer4_node3_MUX_bit_math_h_l1395_c3_68f4_return_output;

     -- layer4_node0_MUX[bit_math_h_l1362_c3_fa41] LATENCY=0
     -- Inputs
     layer4_node0_MUX_bit_math_h_l1362_c3_fa41_cond <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_cond;
     layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iftrue <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iftrue;
     layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iffalse <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_iffalse;
     -- Outputs
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_return_output := layer4_node0_MUX_bit_math_h_l1362_c3_fa41_return_output;

     -- layer4_node1_MUX[bit_math_h_l1373_c3_223f] LATENCY=0
     -- Inputs
     layer4_node1_MUX_bit_math_h_l1373_c3_223f_cond <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_cond;
     layer4_node1_MUX_bit_math_h_l1373_c3_223f_iftrue <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_iftrue;
     layer4_node1_MUX_bit_math_h_l1373_c3_223f_iffalse <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_iffalse;
     -- Outputs
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_return_output := layer4_node1_MUX_bit_math_h_l1373_c3_223f_return_output;

     -- layer4_node2_MUX[bit_math_h_l1384_c3_470b] LATENCY=0
     -- Inputs
     layer4_node2_MUX_bit_math_h_l1384_c3_470b_cond <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_cond;
     layer4_node2_MUX_bit_math_h_l1384_c3_470b_iftrue <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_iftrue;
     layer4_node2_MUX_bit_math_h_l1384_c3_470b_iffalse <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_iffalse;
     -- Outputs
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_return_output := layer4_node2_MUX_bit_math_h_l1384_c3_470b_return_output;

     -- Submodule level 6
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iffalse := VAR_layer4_node0_MUX_bit_math_h_l1362_c3_fa41_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iftrue := VAR_layer4_node1_MUX_bit_math_h_l1373_c3_223f_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iffalse := VAR_layer4_node2_MUX_bit_math_h_l1384_c3_470b_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iftrue := VAR_layer4_node3_MUX_bit_math_h_l1395_c3_68f4_return_output;
     -- layer5_node0_MUX[bit_math_h_l1412_c3_e3bb] LATENCY=0
     -- Inputs
     layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_cond <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_cond;
     layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iftrue <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iftrue;
     layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iffalse <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_iffalse;
     -- Outputs
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_return_output := layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_return_output;

     -- layer5_node1_MUX[bit_math_h_l1423_c3_47e8] LATENCY=0
     -- Inputs
     layer5_node1_MUX_bit_math_h_l1423_c3_47e8_cond <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_cond;
     layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iftrue <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iftrue;
     layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iffalse <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_iffalse;
     -- Outputs
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_return_output := layer5_node1_MUX_bit_math_h_l1423_c3_47e8_return_output;

     -- Submodule level 7
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_iffalse := VAR_layer5_node0_MUX_bit_math_h_l1412_c3_e3bb_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_iftrue := VAR_layer5_node1_MUX_bit_math_h_l1423_c3_47e8_return_output;
     -- layer6_node0_MUX[bit_math_h_l1440_c3_7682] LATENCY=0
     -- Inputs
     layer6_node0_MUX_bit_math_h_l1440_c3_7682_cond <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_cond;
     layer6_node0_MUX_bit_math_h_l1440_c3_7682_iftrue <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_iftrue;
     layer6_node0_MUX_bit_math_h_l1440_c3_7682_iffalse <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_iffalse;
     -- Outputs
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_return_output := layer6_node0_MUX_bit_math_h_l1440_c3_7682_return_output;

     -- Submodule level 8
     VAR_return_output := VAR_layer6_node0_MUX_bit_math_h_l1440_c3_7682_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
