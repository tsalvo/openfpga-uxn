-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 49
entity dei_0CLK_2a8f2cfd is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_device_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dei_0CLK_2a8f2cfd;
architecture arch of dei_0CLK_2a8f2cfd is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal has_written_to_t : unsigned(0 downto 0) := to_unsigned(0, 1);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal device_in_result : device_in_result_t := device_in_result_t_NULL;
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_has_written_to_t : unsigned(0 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_device_in_result : device_in_result_t;
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l408_c6_3838]
signal BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l424_c7_f51a]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l408_c2_ee32]
signal has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l408_c2_ee32]
signal device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : device_in_result_t;

-- t8_MUX[uxn_opcodes_h_l408_c2_ee32]
signal t8_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(3 downto 0);

-- result_is_device_ram_write_MUX[uxn_opcodes_h_l408_c2_ee32]
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
signal result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l424_c11_40d8]
signal BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l427_c1_23a8]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l424_c7_f51a]
signal has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l424_c7_f51a]
signal device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : device_in_result_t;

-- t8_MUX[uxn_opcodes_h_l424_c7_f51a]
signal t8_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l424_c7_f51a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l424_c7_f51a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l424_c7_f51a]
signal result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l424_c7_f51a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l424_c7_f51a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l424_c7_f51a]
signal result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l425_c30_12f3]
signal sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l429_c9_f244]
signal BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l429_c9_ab00]
signal MUX_uxn_opcodes_h_l429_c9_ab00_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l429_c9_ab00_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l429_c9_ab00_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l429_c9_ab00_return_output : unsigned(7 downto 0);

-- UNARY_OP_NOT[uxn_opcodes_h_l430_c8_9d82]
signal UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l430_c1_941a]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l430_c3_b4ff]
signal has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(0 downto 0);

-- device_in_result_MUX[uxn_opcodes_h_l430_c3_b4ff]
signal device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
signal device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : device_in_result_t;
signal device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : device_in_result_t;

-- result_is_opc_done_MUX[uxn_opcodes_h_l430_c3_b4ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l430_c3_b4ff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(0 downto 0);

-- result_device_ram_address_MUX[uxn_opcodes_h_l430_c3_b4ff]
signal result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(7 downto 0);
signal result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l430_c3_b4ff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l430_c3_b4ff]
signal result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(7 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l431_c37_bf4c]
signal BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_right : unsigned(1 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_return_output : unsigned(7 downto 0);

-- device_in[uxn_opcodes_h_l431_c23_7aa9]
signal device_in_uxn_opcodes_h_l431_c23_7aa9_CLOCK_ENABLE : unsigned(0 downto 0);
signal device_in_uxn_opcodes_h_l431_c23_7aa9_device_address : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l431_c23_7aa9_phase : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l431_c23_7aa9_previous_device_ram_read : unsigned(7 downto 0);
signal device_in_uxn_opcodes_h_l431_c23_7aa9_return_output : device_in_result_t;

-- UNARY_OP_NOT[uxn_opcodes_h_l434_c9_825a]
signal UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output : unsigned(0 downto 0);

-- has_written_to_t_MUX[uxn_opcodes_h_l434_c4_9c87]
signal has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(0 downto 0);
signal has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l434_c4_9c87]
signal result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l434_c4_9c87]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l434_c4_9c87]
signal result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l434_c4_9c87]
signal result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(0 downto 0);

function CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6( ref_toks_0 : device_in_result_t;
 ref_toks_1 : unsigned) return device_in_result_t is
 
  variable base : device_in_result_t; 
  variable return_output : device_in_result_t;
begin
      base := ref_toks_0;
      base.is_dei_done := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_bcca( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.device_ram_address := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;
      base.stack_address_sp_offset := ref_toks_10;
      base.is_device_ram_write := ref_toks_11;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838
BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_left,
BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_right,
BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32
has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32
device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- t8_MUX_uxn_opcodes_h_l408_c2_ee32
t8_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
t8_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
t8_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
t8_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32
result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32
result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32
result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32
result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32
result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32
result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32
result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32
result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32
result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond,
result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue,
result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse,
result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8
BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_left,
BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_right,
BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a
has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a
device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- t8_MUX_uxn_opcodes_h_l424_c7_f51a
t8_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
t8_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
t8_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
t8_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a
result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a
result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a
result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a
result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a
result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_cond,
result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l425_c30_12f3
sp_relative_shift_uxn_opcodes_h_l425_c30_12f3 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_ins,
sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_x,
sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_y,
sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244
BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_left,
BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_right,
BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_return_output);

-- MUX_uxn_opcodes_h_l429_c9_ab00
MUX_uxn_opcodes_h_l429_c9_ab00 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l429_c9_ab00_cond,
MUX_uxn_opcodes_h_l429_c9_ab00_iftrue,
MUX_uxn_opcodes_h_l429_c9_ab00_iffalse,
MUX_uxn_opcodes_h_l429_c9_ab00_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82
UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_expr,
UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff
has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_cond,
has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output);

-- device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff
device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff : entity work.MUX_uint1_t_device_in_result_t_device_in_result_t_0CLK_de264c78 port map (
device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_cond,
device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue,
device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse,
device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff
result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff
result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output);

-- result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff
result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_cond,
result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue,
result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse,
result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff
result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_cond,
result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c
BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c : entity work.BIN_OP_MINUS_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_left,
BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_right,
BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_return_output);

-- device_in_uxn_opcodes_h_l431_c23_7aa9
device_in_uxn_opcodes_h_l431_c23_7aa9 : entity work.device_in_0CLK_85463cfa port map (
clk,
device_in_uxn_opcodes_h_l431_c23_7aa9_CLOCK_ENABLE,
device_in_uxn_opcodes_h_l431_c23_7aa9_device_address,
device_in_uxn_opcodes_h_l431_c23_7aa9_phase,
device_in_uxn_opcodes_h_l431_c23_7aa9_previous_device_ram_read,
device_in_uxn_opcodes_h_l431_c23_7aa9_return_output);

-- UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a
UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_expr,
UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output);

-- has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87
has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_cond,
has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue,
has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse,
has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87
result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_cond,
result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87
result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87
result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_device_ram_read,
 -- Registers
 has_written_to_t,
 t8,
 device_in_result,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 t8_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 t8_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_return_output,
 sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_return_output,
 MUX_uxn_opcodes_h_l429_c9_ab00_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output,
 device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output,
 result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_return_output,
 device_in_uxn_opcodes_h_l431_c23_7aa9_return_output,
 UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output,
 has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : device_in_result_t;
 variable VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l408_c2_ee32_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l413_c3_a0fb : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l419_c3_4291 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output : unsigned(0 downto 0);
 variable VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l428_c3_c09b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l429_c9_ab00_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l429_c9_ab00_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l429_c9_ab00_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l429_c9_ab00_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l430_c8_0c2d_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : device_in_result_t;
 variable VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_cond : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_device_address : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_phase : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_previous_device_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_return_output : unsigned(7 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_return_output : device_in_result_t;
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l432_c32_858a_return_output : unsigned(7 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(0 downto 0);
 variable VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l436_c5_7a3b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l437_c23_80bd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l430_l408_l424_DUPLICATE_35e2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l430_l408_l434_l424_DUPLICATE_2ecd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2873_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l430_l424_DUPLICATE_21df_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2594_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_bcca_uxn_opcodes_h_l446_l402_DUPLICATE_432a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_has_written_to_t : unsigned(0 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_device_in_result : device_in_result_t;
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_has_written_to_t := has_written_to_t;
  REG_VAR_t8 := t8;
  REG_VAR_device_in_result := device_in_result;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iffalse := to_unsigned(0, 1);
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l436_c5_7a3b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l436_c5_7a3b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := to_unsigned(0, 1);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_right := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l419_c3_4291 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l419_c3_4291;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_right := to_unsigned(2, 2);
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l428_c3_c09b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_result_sp_relative_shift_uxn_opcodes_h_l428_c3_c09b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l413_c3_a0fb := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l413_c3_a0fb;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_device_ram_read := previous_device_ram_read;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_CLOCK_ENABLE;
     VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := device_in_result;
     VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse := device_in_result;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_expr := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue := has_written_to_t;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse := has_written_to_t;
     VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_left := VAR_phase;
     VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_previous_device_ram_read := VAR_previous_device_ram_read;
     VAR_MUX_uxn_opcodes_h_l429_c9_ab00_iftrue := VAR_previous_stack_read;
     VAR_MUX_uxn_opcodes_h_l429_c9_ab00_iffalse := t8;
     VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := t8;
     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l424_c11_40d8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_left;
     BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output := BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l430_l408_l424_DUPLICATE_35e2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l430_l408_l424_DUPLICATE_35e2_return_output := result.device_ram_address;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l408_c2_ee32_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l408_c2_ee32_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d[uxn_opcodes_h_l437_c23_80bd] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l437_c23_80bd_return_output := device_in_result.dei_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2873 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2873_return_output := result.is_opc_done;

     -- BIN_OP_MINUS[uxn_opcodes_h_l431_c37_bf4c] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_left;
     BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_return_output := BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l408_c6_3838] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_left;
     BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output := BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l430_l408_l434_l424_DUPLICATE_2ecd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l430_l408_l434_l424_DUPLICATE_2ecd_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l425_c30_12f3] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_ins;
     sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_x <= VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_x;
     sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_y <= VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_return_output := sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_return_output;

     -- result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output := result.is_device_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d[uxn_opcodes_h_l430_c8_0c2d] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l430_c8_0c2d_return_output := device_in_result.is_dei_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2594 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2594_return_output := result.stack_address_sp_offset;

     -- UNARY_OP_NOT[uxn_opcodes_h_l434_c9_825a] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output := UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l430_l424_DUPLICATE_21df LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l430_l424_DUPLICATE_21df_return_output := result.is_stack_write;

     -- device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l408_c2_ee32_return_output := CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6(
     device_in_result,
     to_unsigned(0, 1));

     -- BIN_OP_EQ[uxn_opcodes_h_l429_c9_f244] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_left;
     BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_return_output := BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l408_c6_3838_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l424_c11_40d8_return_output;
     VAR_MUX_uxn_opcodes_h_l429_c9_ab00_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l429_c9_f244_return_output;
     VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_phase := VAR_BIN_OP_MINUS_uxn_opcodes_h_l431_c37_bf4c_return_output;
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_expr := VAR_CONST_REF_RD_uint1_t_device_in_result_t_is_dei_done_d41d_uxn_opcodes_h_l430_c8_0c2d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2873_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2873_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2873_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l430_l424_DUPLICATE_21df_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l430_l424_DUPLICATE_21df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2594_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2594_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l430_l434_l424_DUPLICATE_2594_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_dei_value_d41d_uxn_opcodes_h_l437_c23_80bd_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l430_l408_l424_DUPLICATE_35e2_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l430_l408_l424_DUPLICATE_35e2_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_device_ram_address_d41d_uxn_opcodes_h_l430_l408_l424_DUPLICATE_35e2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l430_l408_l434_l424_DUPLICATE_2ecd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l430_l408_l434_l424_DUPLICATE_2ecd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l430_l408_l434_l424_DUPLICATE_2ecd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l430_l408_l434_l424_DUPLICATE_2ecd_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l434_c9_825a_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue := VAR_device_in_result_TRUE_INPUT_MUX_CONST_REF_RD_device_in_result_t_device_in_result_t_6bb6_uxn_opcodes_h_l408_c2_ee32_return_output;
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_is_device_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_device_ram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l408_c2_ee32_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l408_c2_ee32_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l408_c2_ee32_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l425_c30_12f3_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l434_c4_9c87] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_return_output := has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;

     -- UNARY_OP_NOT[uxn_opcodes_h_l430_c8_9d82] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_expr <= VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output := UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- MUX[uxn_opcodes_h_l429_c9_ab00] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l429_c9_ab00_cond <= VAR_MUX_uxn_opcodes_h_l429_c9_ab00_cond;
     MUX_uxn_opcodes_h_l429_c9_ab00_iftrue <= VAR_MUX_uxn_opcodes_h_l429_c9_ab00_iftrue;
     MUX_uxn_opcodes_h_l429_c9_ab00_iffalse <= VAR_MUX_uxn_opcodes_h_l429_c9_ab00_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l429_c9_ab00_return_output := MUX_uxn_opcodes_h_l429_c9_ab00_return_output;

     -- result_is_device_ram_write_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l434_c4_9c87] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l434_c4_9c87] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l434_c4_9c87] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l434_c4_9c87] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_cond;
     result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_return_output := result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_device_address := VAR_MUX_uxn_opcodes_h_l429_c9_ab00_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_MUX_uxn_opcodes_h_l429_c9_ab00_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_cond := VAR_UNARY_OP_NOT_uxn_opcodes_h_l430_c8_9d82_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l434_c4_9c87_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l430_c3_b4ff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l430_c3_b4ff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output := result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l430_c3_b4ff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l430_c3_b4ff] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output := has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l430_c3_b4ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l427_c1_23a8] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_return_output;

     -- t8_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     t8_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     t8_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := t8_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l427_c1_23a8_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_t8_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- has_written_to_t_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- t8_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     t8_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     t8_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := t8_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l430_c1_941a] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_return_output;

     -- Submodule level 4
     VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l430_c1_941a_return_output;
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_has_written_to_t_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;
     -- has_written_to_t_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- device_in[uxn_opcodes_h_l431_c23_7aa9] LATENCY=0
     -- Clock enable
     device_in_uxn_opcodes_h_l431_c23_7aa9_CLOCK_ENABLE <= VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_CLOCK_ENABLE;
     -- Inputs
     device_in_uxn_opcodes_h_l431_c23_7aa9_device_address <= VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_device_address;
     device_in_uxn_opcodes_h_l431_c23_7aa9_phase <= VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_phase;
     device_in_uxn_opcodes_h_l431_c23_7aa9_previous_device_ram_read <= VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_previous_device_ram_read;
     -- Outputs
     VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_return_output := device_in_uxn_opcodes_h_l431_c23_7aa9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- Submodule level 5
     VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue := VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_return_output;
     REG_VAR_has_written_to_t := VAR_has_written_to_t_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l430_c3_b4ff] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_cond;
     device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output := device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;

     -- CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d[uxn_opcodes_h_l432_c32_858a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l432_c32_858a_return_output := VAR_device_in_uxn_opcodes_h_l431_c23_7aa9_return_output.device_ram_address;

     -- Submodule level 6
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue := VAR_CONST_REF_RD_uint8_t_device_in_result_t_device_ram_address_d41d_uxn_opcodes_h_l432_c32_858a_return_output;
     VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l430_c3_b4ff] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;

     -- device_in_result_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- Submodule level 7
     VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_device_in_result_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l430_c3_b4ff_return_output;
     -- device_in_result_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- result_device_ram_address_MUX[uxn_opcodes_h_l424_c7_f51a] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;

     -- Submodule level 8
     REG_VAR_device_in_result := VAR_device_in_result_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse := VAR_result_device_ram_address_MUX_uxn_opcodes_h_l424_c7_f51a_return_output;
     -- result_device_ram_address_MUX[uxn_opcodes_h_l408_c2_ee32] LATENCY=0
     -- Inputs
     result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_cond <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_cond;
     result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iftrue;
     result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse <= VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_iffalse;
     -- Outputs
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_return_output := result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_bcca_uxn_opcodes_h_l446_l402_DUPLICATE_432a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_bcca_uxn_opcodes_h_l446_l402_DUPLICATE_432a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_bcca(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_device_ram_address_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l408_c2_ee32_return_output,
     VAR_result_is_device_ram_write_MUX_uxn_opcodes_h_l408_c2_ee32_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_bcca_uxn_opcodes_h_l446_l402_DUPLICATE_432a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_bcca_uxn_opcodes_h_l446_l402_DUPLICATE_432a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_has_written_to_t <= REG_VAR_has_written_to_t;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_device_in_result <= REG_VAR_device_in_result;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     has_written_to_t <= REG_COMB_has_written_to_t;
     t8 <= REG_COMB_t8;
     device_in_result <= REG_COMB_device_in_result;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
