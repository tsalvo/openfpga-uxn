-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity lth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_226c8821;
architecture arch of lth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1912_c6_fef5]
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1912_c2_5073]
signal t8_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1912_c2_5073]
signal n8_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1912_c2_5073]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1925_c11_ffe9]
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1925_c7_c37b]
signal t8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1925_c7_c37b]
signal n8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1925_c7_c37b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1925_c7_c37b]
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1925_c7_c37b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1925_c7_c37b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1925_c7_c37b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1928_c11_8292]
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1928_c7_a9fc]
signal t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1928_c7_a9fc]
signal n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1928_c7_a9fc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1928_c7_a9fc]
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1928_c7_a9fc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1928_c7_a9fc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1928_c7_a9fc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1931_c11_d814]
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1931_c7_a5e3]
signal n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1931_c7_a5e3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1931_c7_a5e3]
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1931_c7_a5e3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1931_c7_a5e3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1931_c7_a5e3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1933_c30_d240]
signal sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1936_c21_b109]
signal BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1936_c21_3c13]
signal MUX_uxn_opcodes_h_l1936_c21_3c13_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1936_c21_3c13_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1936_c21_3c13_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1936_c21_3c13_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5
BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_left,
BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_right,
BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output);

-- t8_MUX_uxn_opcodes_h_l1912_c2_5073
t8_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
t8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
t8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
t8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- n8_MUX_uxn_opcodes_h_l1912_c2_5073
n8_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
n8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
n8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
n8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_left,
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_right,
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output);

-- t8_MUX_uxn_opcodes_h_l1925_c7_c37b
t8_MUX_uxn_opcodes_h_l1925_c7_c37b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond,
t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue,
t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse,
t8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output);

-- n8_MUX_uxn_opcodes_h_l1925_c7_c37b
n8_MUX_uxn_opcodes_h_l1925_c7_c37b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond,
n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue,
n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse,
n8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_left,
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_right,
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output);

-- t8_MUX_uxn_opcodes_h_l1928_c7_a9fc
t8_MUX_uxn_opcodes_h_l1928_c7_a9fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond,
t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue,
t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse,
t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output);

-- n8_MUX_uxn_opcodes_h_l1928_c7_a9fc
n8_MUX_uxn_opcodes_h_l1928_c7_a9fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond,
n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue,
n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse,
n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_left,
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_right,
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output);

-- n8_MUX_uxn_opcodes_h_l1931_c7_a5e3
n8_MUX_uxn_opcodes_h_l1931_c7_a5e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond,
n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue,
n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse,
n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1933_c30_d240
sp_relative_shift_uxn_opcodes_h_l1933_c30_d240 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_ins,
sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_x,
sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_y,
sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109
BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_left,
BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_right,
BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_return_output);

-- MUX_uxn_opcodes_h_l1936_c21_3c13
MUX_uxn_opcodes_h_l1936_c21_3c13 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1936_c21_3c13_cond,
MUX_uxn_opcodes_h_l1936_c21_3c13_iftrue,
MUX_uxn_opcodes_h_l1936_c21_3c13_iffalse,
MUX_uxn_opcodes_h_l1936_c21_3c13_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output,
 t8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 n8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output,
 t8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output,
 n8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output,
 t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output,
 n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output,
 n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output,
 sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_return_output,
 MUX_uxn_opcodes_h_l1936_c21_3c13_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1917_c3_a587 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_6e92 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_88d2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1935_c3_4e34 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1912_l1931_l1925_l1928_DUPLICATE_de19_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_92b6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_9401_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_2dd0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1931_l1928_DUPLICATE_7da1_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1940_l1908_DUPLICATE_69d5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_88d2 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_88d2;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_6e92 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_6e92;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1935_c3_4e34 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1935_c3_4e34;
     VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1917_c3_a587 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1917_c3_a587;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse := t8;
     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1912_c2_5073_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_9401 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_9401_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1931_c11_d814] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_left;
     BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output := BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1912_l1931_l1925_l1928_DUPLICATE_de19 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1912_l1931_l1925_l1928_DUPLICATE_de19_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l1933_c30_d240] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_ins;
     sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_x;
     sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_return_output := sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1912_c2_5073_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1931_l1928_DUPLICATE_7da1 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1931_l1928_DUPLICATE_7da1_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1925_c11_ffe9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1912_c2_5073_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_92b6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_92b6_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1912_c2_5073_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1928_c11_8292] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_left;
     BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output := BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1912_c6_fef5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_2dd0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_2dd0_return_output := result.is_stack_write;

     -- BIN_OP_LT[uxn_opcodes_h_l1936_c21_b109] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_left;
     BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_return_output := BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1912_c6_fef5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_ffe9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8292_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_d814_return_output;
     VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1936_c21_b109_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_9401_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_9401_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_9401_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_92b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_92b6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_92b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_2dd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_2dd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1931_l1925_l1928_DUPLICATE_2dd0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1931_l1928_DUPLICATE_7da1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1931_l1928_DUPLICATE_7da1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1912_l1931_l1925_l1928_DUPLICATE_de19_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1912_l1931_l1925_l1928_DUPLICATE_de19_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1912_l1931_l1925_l1928_DUPLICATE_de19_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1912_l1931_l1925_l1928_DUPLICATE_de19_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1912_c2_5073_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1912_c2_5073_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1912_c2_5073_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1912_c2_5073_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1933_c30_d240_return_output;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1931_c7_a5e3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1931_c7_a5e3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1931_c7_a5e3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;

     -- MUX[uxn_opcodes_h_l1936_c21_3c13] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1936_c21_3c13_cond <= VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_cond;
     MUX_uxn_opcodes_h_l1936_c21_3c13_iftrue <= VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_iftrue;
     MUX_uxn_opcodes_h_l1936_c21_3c13_iffalse <= VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_return_output := MUX_uxn_opcodes_h_l1936_c21_3c13_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1931_c7_a5e3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1931_c7_a5e3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond;
     n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue;
     n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output := n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1928_c7_a9fc] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond <= VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond;
     t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue;
     t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output := t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue := VAR_MUX_uxn_opcodes_h_l1936_c21_3c13_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1931_c7_a5e3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1928_c7_a9fc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;

     -- n8_MUX[uxn_opcodes_h_l1928_c7_a9fc] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond;
     n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue;
     n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output := n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1928_c7_a9fc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1928_c7_a9fc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;

     -- t8_MUX[uxn_opcodes_h_l1925_c7_c37b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond;
     t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue;
     t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output := t8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1928_c7_a9fc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_a5e3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;
     -- n8_MUX[uxn_opcodes_h_l1925_c7_c37b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_cond;
     n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue;
     n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output := n8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     t8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     t8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := t8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1925_c7_c37b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1925_c7_c37b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1925_c7_c37b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1928_c7_a9fc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output := result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1925_c7_c37b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_a9fc_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1925_c7_c37b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- n8_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     n8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     n8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := n8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_c37b_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1912_c2_5073] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_return_output := result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1940_l1908_DUPLICATE_69d5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1940_l1908_DUPLICATE_69d5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1912_c2_5073_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1912_c2_5073_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1940_l1908_DUPLICATE_69d5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1940_l1908_DUPLICATE_69d5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
