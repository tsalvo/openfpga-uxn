-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_226c8821;
architecture arch of equ_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1163_c6_07fa]
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal n8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal t8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1163_c2_5c09]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1176_c11_8a1d]
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1176_c7_f17a]
signal n8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1176_c7_f17a]
signal t8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1176_c7_f17a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1176_c7_f17a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1176_c7_f17a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1176_c7_f17a]
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1176_c7_f17a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1179_c11_5041]
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1179_c7_a9f9]
signal n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1179_c7_a9f9]
signal t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1179_c7_a9f9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1179_c7_a9f9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1179_c7_a9f9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1179_c7_a9f9]
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1179_c7_a9f9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1182_c11_4a85]
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1182_c7_f007]
signal n8_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1182_c7_f007]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1182_c7_f007]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1182_c7_f007]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1182_c7_f007]
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1182_c7_f007]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1184_c30_4e3b]
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1187_c21_9362]
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1187_c21_43ae]
signal MUX_uxn_opcodes_h_l1187_c21_43ae_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_43ae_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_43ae_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1187_c21_43ae_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a6df( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_left,
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_right,
BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output);

-- n8_MUX_uxn_opcodes_h_l1163_c2_5c09
n8_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
n8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- t8_MUX_uxn_opcodes_h_l1163_c2_5c09
t8_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
t8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_left,
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_right,
BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output);

-- n8_MUX_uxn_opcodes_h_l1176_c7_f17a
n8_MUX_uxn_opcodes_h_l1176_c7_f17a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond,
n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue,
n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse,
n8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output);

-- t8_MUX_uxn_opcodes_h_l1176_c7_f17a
t8_MUX_uxn_opcodes_h_l1176_c7_f17a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond,
t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue,
t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse,
t8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_left,
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_right,
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output);

-- n8_MUX_uxn_opcodes_h_l1179_c7_a9f9
n8_MUX_uxn_opcodes_h_l1179_c7_a9f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond,
n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue,
n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse,
n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output);

-- t8_MUX_uxn_opcodes_h_l1179_c7_a9f9
t8_MUX_uxn_opcodes_h_l1179_c7_a9f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond,
t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue,
t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse,
t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_left,
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_right,
BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output);

-- n8_MUX_uxn_opcodes_h_l1182_c7_f007
n8_MUX_uxn_opcodes_h_l1182_c7_f007 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1182_c7_f007_cond,
n8_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue,
n8_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse,
n8_MUX_uxn_opcodes_h_l1182_c7_f007_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_cond,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b
sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_ins,
sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_x,
sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_y,
sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_left,
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_right,
BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_return_output);

-- MUX_uxn_opcodes_h_l1187_c21_43ae
MUX_uxn_opcodes_h_l1187_c21_43ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1187_c21_43ae_cond,
MUX_uxn_opcodes_h_l1187_c21_43ae_iftrue,
MUX_uxn_opcodes_h_l1187_c21_43ae_iffalse,
MUX_uxn_opcodes_h_l1187_c21_43ae_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output,
 n8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 t8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output,
 n8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output,
 t8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output,
 n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output,
 t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output,
 n8_MUX_uxn_opcodes_h_l1182_c7_f007_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_return_output,
 sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_return_output,
 MUX_uxn_opcodes_h_l1187_c21_43ae_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_b493 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_5f5a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_015f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_5c2a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1179_l1163_l1182_l1176_DUPLICATE_37ec_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_9db0_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_91e1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_0181_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1179_l1182_DUPLICATE_2367_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1159_l1191_DUPLICATE_6eba_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_015f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1177_c3_015f;
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_5f5a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1173_c3_5f5a;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_b493 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1168_c3_b493;
     VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_5c2a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1186_c3_5c2a;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_y := resize(to_signed(-1, 2), 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1187_c21_9362] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_left;
     BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_return_output := BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1179_l1182_DUPLICATE_2367 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1179_l1182_DUPLICATE_2367_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_9db0 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_9db0_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1163_c6_07fa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_left;
     BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output := BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_91e1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_91e1_return_output := result.is_opc_done;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1182_c11_4a85] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_left;
     BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output := BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1176_c11_8a1d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_0181 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_0181_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1179_c11_5041] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_left;
     BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output := BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1179_l1163_l1182_l1176_DUPLICATE_37ec LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1179_l1163_l1182_l1176_DUPLICATE_37ec_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l1184_c30_4e3b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_ins;
     sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_x;
     sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_return_output := sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1163_c6_07fa_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1176_c11_8a1d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_5041_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1182_c11_4a85_return_output;
     VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1187_c21_9362_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_9db0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_9db0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_9db0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_91e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_91e1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_91e1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_0181_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_0181_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1179_l1182_l1176_DUPLICATE_0181_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1179_l1182_DUPLICATE_2367_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1179_l1182_DUPLICATE_2367_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1179_l1163_l1182_l1176_DUPLICATE_37ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1179_l1163_l1182_l1176_DUPLICATE_37ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1179_l1163_l1182_l1176_DUPLICATE_37ec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1179_l1163_l1182_l1176_DUPLICATE_37ec_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1163_c2_5c09_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1184_c30_4e3b_return_output;
     -- MUX[uxn_opcodes_h_l1187_c21_43ae] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1187_c21_43ae_cond <= VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_cond;
     MUX_uxn_opcodes_h_l1187_c21_43ae_iftrue <= VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_iftrue;
     MUX_uxn_opcodes_h_l1187_c21_43ae_iffalse <= VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_return_output := MUX_uxn_opcodes_h_l1187_c21_43ae_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1182_c7_f007] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1182_c7_f007] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1182_c7_f007] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;

     -- t8_MUX[uxn_opcodes_h_l1179_c7_a9f9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond;
     t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue;
     t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output := t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1182_c7_f007] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;

     -- n8_MUX[uxn_opcodes_h_l1182_c7_f007] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1182_c7_f007_cond <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_cond;
     n8_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue;
     n8_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_return_output := n8_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue := VAR_MUX_uxn_opcodes_h_l1187_c21_43ae_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;
     -- n8_MUX[uxn_opcodes_h_l1179_c7_a9f9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond;
     n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue;
     n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output := n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1182_c7_f007] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_return_output := result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1179_c7_a9f9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1176_c7_f17a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond;
     t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue;
     t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output := t8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1179_c7_a9f9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1179_c7_a9f9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1179_c7_a9f9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1182_c7_f007_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1176_c7_f17a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1176_c7_f17a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;

     -- t8_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := t8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1176_c7_f17a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1176_c7_f17a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_cond;
     n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue;
     n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output := n8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1176_c7_f17a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1179_c7_a9f9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_a9f9_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1176_c7_f17a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- n8_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := n8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1176_c7_f17a_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1163_c2_5c09] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output := result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1159_l1191_DUPLICATE_6eba LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1159_l1191_DUPLICATE_6eba_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a6df(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1163_c2_5c09_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1159_l1191_DUPLICATE_6eba_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l1159_l1191_DUPLICATE_6eba_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
