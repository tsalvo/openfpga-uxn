-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 134
entity uint8_mux128_0CLK_9347d63d is
port(
 sel : in unsigned(6 downto 0);
 in0 : in unsigned(7 downto 0);
 in1 : in unsigned(7 downto 0);
 in2 : in unsigned(7 downto 0);
 in3 : in unsigned(7 downto 0);
 in4 : in unsigned(7 downto 0);
 in5 : in unsigned(7 downto 0);
 in6 : in unsigned(7 downto 0);
 in7 : in unsigned(7 downto 0);
 in8 : in unsigned(7 downto 0);
 in9 : in unsigned(7 downto 0);
 in10 : in unsigned(7 downto 0);
 in11 : in unsigned(7 downto 0);
 in12 : in unsigned(7 downto 0);
 in13 : in unsigned(7 downto 0);
 in14 : in unsigned(7 downto 0);
 in15 : in unsigned(7 downto 0);
 in16 : in unsigned(7 downto 0);
 in17 : in unsigned(7 downto 0);
 in18 : in unsigned(7 downto 0);
 in19 : in unsigned(7 downto 0);
 in20 : in unsigned(7 downto 0);
 in21 : in unsigned(7 downto 0);
 in22 : in unsigned(7 downto 0);
 in23 : in unsigned(7 downto 0);
 in24 : in unsigned(7 downto 0);
 in25 : in unsigned(7 downto 0);
 in26 : in unsigned(7 downto 0);
 in27 : in unsigned(7 downto 0);
 in28 : in unsigned(7 downto 0);
 in29 : in unsigned(7 downto 0);
 in30 : in unsigned(7 downto 0);
 in31 : in unsigned(7 downto 0);
 in32 : in unsigned(7 downto 0);
 in33 : in unsigned(7 downto 0);
 in34 : in unsigned(7 downto 0);
 in35 : in unsigned(7 downto 0);
 in36 : in unsigned(7 downto 0);
 in37 : in unsigned(7 downto 0);
 in38 : in unsigned(7 downto 0);
 in39 : in unsigned(7 downto 0);
 in40 : in unsigned(7 downto 0);
 in41 : in unsigned(7 downto 0);
 in42 : in unsigned(7 downto 0);
 in43 : in unsigned(7 downto 0);
 in44 : in unsigned(7 downto 0);
 in45 : in unsigned(7 downto 0);
 in46 : in unsigned(7 downto 0);
 in47 : in unsigned(7 downto 0);
 in48 : in unsigned(7 downto 0);
 in49 : in unsigned(7 downto 0);
 in50 : in unsigned(7 downto 0);
 in51 : in unsigned(7 downto 0);
 in52 : in unsigned(7 downto 0);
 in53 : in unsigned(7 downto 0);
 in54 : in unsigned(7 downto 0);
 in55 : in unsigned(7 downto 0);
 in56 : in unsigned(7 downto 0);
 in57 : in unsigned(7 downto 0);
 in58 : in unsigned(7 downto 0);
 in59 : in unsigned(7 downto 0);
 in60 : in unsigned(7 downto 0);
 in61 : in unsigned(7 downto 0);
 in62 : in unsigned(7 downto 0);
 in63 : in unsigned(7 downto 0);
 in64 : in unsigned(7 downto 0);
 in65 : in unsigned(7 downto 0);
 in66 : in unsigned(7 downto 0);
 in67 : in unsigned(7 downto 0);
 in68 : in unsigned(7 downto 0);
 in69 : in unsigned(7 downto 0);
 in70 : in unsigned(7 downto 0);
 in71 : in unsigned(7 downto 0);
 in72 : in unsigned(7 downto 0);
 in73 : in unsigned(7 downto 0);
 in74 : in unsigned(7 downto 0);
 in75 : in unsigned(7 downto 0);
 in76 : in unsigned(7 downto 0);
 in77 : in unsigned(7 downto 0);
 in78 : in unsigned(7 downto 0);
 in79 : in unsigned(7 downto 0);
 in80 : in unsigned(7 downto 0);
 in81 : in unsigned(7 downto 0);
 in82 : in unsigned(7 downto 0);
 in83 : in unsigned(7 downto 0);
 in84 : in unsigned(7 downto 0);
 in85 : in unsigned(7 downto 0);
 in86 : in unsigned(7 downto 0);
 in87 : in unsigned(7 downto 0);
 in88 : in unsigned(7 downto 0);
 in89 : in unsigned(7 downto 0);
 in90 : in unsigned(7 downto 0);
 in91 : in unsigned(7 downto 0);
 in92 : in unsigned(7 downto 0);
 in93 : in unsigned(7 downto 0);
 in94 : in unsigned(7 downto 0);
 in95 : in unsigned(7 downto 0);
 in96 : in unsigned(7 downto 0);
 in97 : in unsigned(7 downto 0);
 in98 : in unsigned(7 downto 0);
 in99 : in unsigned(7 downto 0);
 in100 : in unsigned(7 downto 0);
 in101 : in unsigned(7 downto 0);
 in102 : in unsigned(7 downto 0);
 in103 : in unsigned(7 downto 0);
 in104 : in unsigned(7 downto 0);
 in105 : in unsigned(7 downto 0);
 in106 : in unsigned(7 downto 0);
 in107 : in unsigned(7 downto 0);
 in108 : in unsigned(7 downto 0);
 in109 : in unsigned(7 downto 0);
 in110 : in unsigned(7 downto 0);
 in111 : in unsigned(7 downto 0);
 in112 : in unsigned(7 downto 0);
 in113 : in unsigned(7 downto 0);
 in114 : in unsigned(7 downto 0);
 in115 : in unsigned(7 downto 0);
 in116 : in unsigned(7 downto 0);
 in117 : in unsigned(7 downto 0);
 in118 : in unsigned(7 downto 0);
 in119 : in unsigned(7 downto 0);
 in120 : in unsigned(7 downto 0);
 in121 : in unsigned(7 downto 0);
 in122 : in unsigned(7 downto 0);
 in123 : in unsigned(7 downto 0);
 in124 : in unsigned(7 downto 0);
 in125 : in unsigned(7 downto 0);
 in126 : in unsigned(7 downto 0);
 in127 : in unsigned(7 downto 0);
 return_output : out unsigned(7 downto 0));
end uint8_mux128_0CLK_9347d63d;
architecture arch of uint8_mux128_0CLK_9347d63d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_8bd4]
signal layer0_node0_MUX_bit_math_h_l18_c3_8bd4_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iftrue : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iffalse : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_8bd4_return_output : unsigned(7 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_b2fc]
signal layer0_node1_MUX_bit_math_h_l29_c3_b2fc_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iftrue : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iffalse : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_b2fc_return_output : unsigned(7 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_3d12]
signal layer0_node2_MUX_bit_math_h_l40_c3_3d12_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_3d12_iftrue : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_3d12_iffalse : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_3d12_return_output : unsigned(7 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_13b9]
signal layer0_node3_MUX_bit_math_h_l51_c3_13b9_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_13b9_iftrue : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_13b9_iffalse : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_13b9_return_output : unsigned(7 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_be4c]
signal layer0_node4_MUX_bit_math_h_l62_c3_be4c_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_be4c_iftrue : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_be4c_iffalse : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_be4c_return_output : unsigned(7 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_936b]
signal layer0_node5_MUX_bit_math_h_l73_c3_936b_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_936b_iftrue : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_936b_iffalse : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_936b_return_output : unsigned(7 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_6f9a]
signal layer0_node6_MUX_bit_math_h_l84_c3_6f9a_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iftrue : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iffalse : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_6f9a_return_output : unsigned(7 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_f259]
signal layer0_node7_MUX_bit_math_h_l95_c3_f259_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_f259_iftrue : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_f259_iffalse : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_f259_return_output : unsigned(7 downto 0);

-- layer0_node8_MUX[bit_math_h_l106_c3_2e0c]
signal layer0_node8_MUX_bit_math_h_l106_c3_2e0c_cond : unsigned(0 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iftrue : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iffalse : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_2e0c_return_output : unsigned(7 downto 0);

-- layer0_node9_MUX[bit_math_h_l117_c3_1a47]
signal layer0_node9_MUX_bit_math_h_l117_c3_1a47_cond : unsigned(0 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_1a47_iftrue : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_1a47_iffalse : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_1a47_return_output : unsigned(7 downto 0);

-- layer0_node10_MUX[bit_math_h_l128_c3_0e40]
signal layer0_node10_MUX_bit_math_h_l128_c3_0e40_cond : unsigned(0 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_0e40_iftrue : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_0e40_iffalse : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_0e40_return_output : unsigned(7 downto 0);

-- layer0_node11_MUX[bit_math_h_l139_c3_381c]
signal layer0_node11_MUX_bit_math_h_l139_c3_381c_cond : unsigned(0 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_381c_iftrue : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_381c_iffalse : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_381c_return_output : unsigned(7 downto 0);

-- layer0_node12_MUX[bit_math_h_l150_c3_1560]
signal layer0_node12_MUX_bit_math_h_l150_c3_1560_cond : unsigned(0 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_1560_iftrue : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_1560_iffalse : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_1560_return_output : unsigned(7 downto 0);

-- layer0_node13_MUX[bit_math_h_l161_c3_3a1c]
signal layer0_node13_MUX_bit_math_h_l161_c3_3a1c_cond : unsigned(0 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iftrue : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iffalse : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_3a1c_return_output : unsigned(7 downto 0);

-- layer0_node14_MUX[bit_math_h_l172_c3_7ef7]
signal layer0_node14_MUX_bit_math_h_l172_c3_7ef7_cond : unsigned(0 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iftrue : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iffalse : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_7ef7_return_output : unsigned(7 downto 0);

-- layer0_node15_MUX[bit_math_h_l183_c3_392b]
signal layer0_node15_MUX_bit_math_h_l183_c3_392b_cond : unsigned(0 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_392b_iftrue : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_392b_iffalse : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_392b_return_output : unsigned(7 downto 0);

-- layer0_node16_MUX[bit_math_h_l194_c3_cada]
signal layer0_node16_MUX_bit_math_h_l194_c3_cada_cond : unsigned(0 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_cada_iftrue : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_cada_iffalse : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_cada_return_output : unsigned(7 downto 0);

-- layer0_node17_MUX[bit_math_h_l205_c3_39fd]
signal layer0_node17_MUX_bit_math_h_l205_c3_39fd_cond : unsigned(0 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_39fd_iftrue : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_39fd_iffalse : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_39fd_return_output : unsigned(7 downto 0);

-- layer0_node18_MUX[bit_math_h_l216_c3_23c8]
signal layer0_node18_MUX_bit_math_h_l216_c3_23c8_cond : unsigned(0 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_23c8_iftrue : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_23c8_iffalse : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_23c8_return_output : unsigned(7 downto 0);

-- layer0_node19_MUX[bit_math_h_l227_c3_ea58]
signal layer0_node19_MUX_bit_math_h_l227_c3_ea58_cond : unsigned(0 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_ea58_iftrue : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_ea58_iffalse : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_ea58_return_output : unsigned(7 downto 0);

-- layer0_node20_MUX[bit_math_h_l238_c3_eb78]
signal layer0_node20_MUX_bit_math_h_l238_c3_eb78_cond : unsigned(0 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_eb78_iftrue : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_eb78_iffalse : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_eb78_return_output : unsigned(7 downto 0);

-- layer0_node21_MUX[bit_math_h_l249_c3_228d]
signal layer0_node21_MUX_bit_math_h_l249_c3_228d_cond : unsigned(0 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_228d_iftrue : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_228d_iffalse : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_228d_return_output : unsigned(7 downto 0);

-- layer0_node22_MUX[bit_math_h_l260_c3_1c3c]
signal layer0_node22_MUX_bit_math_h_l260_c3_1c3c_cond : unsigned(0 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iftrue : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iffalse : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_1c3c_return_output : unsigned(7 downto 0);

-- layer0_node23_MUX[bit_math_h_l271_c3_6340]
signal layer0_node23_MUX_bit_math_h_l271_c3_6340_cond : unsigned(0 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_6340_iftrue : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_6340_iffalse : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_6340_return_output : unsigned(7 downto 0);

-- layer0_node24_MUX[bit_math_h_l282_c3_670b]
signal layer0_node24_MUX_bit_math_h_l282_c3_670b_cond : unsigned(0 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_670b_iftrue : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_670b_iffalse : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_670b_return_output : unsigned(7 downto 0);

-- layer0_node25_MUX[bit_math_h_l293_c3_83e8]
signal layer0_node25_MUX_bit_math_h_l293_c3_83e8_cond : unsigned(0 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_83e8_iftrue : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_83e8_iffalse : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_83e8_return_output : unsigned(7 downto 0);

-- layer0_node26_MUX[bit_math_h_l304_c3_53e2]
signal layer0_node26_MUX_bit_math_h_l304_c3_53e2_cond : unsigned(0 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_53e2_iftrue : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_53e2_iffalse : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_53e2_return_output : unsigned(7 downto 0);

-- layer0_node27_MUX[bit_math_h_l315_c3_ac24]
signal layer0_node27_MUX_bit_math_h_l315_c3_ac24_cond : unsigned(0 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_ac24_iftrue : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_ac24_iffalse : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_ac24_return_output : unsigned(7 downto 0);

-- layer0_node28_MUX[bit_math_h_l326_c3_97ed]
signal layer0_node28_MUX_bit_math_h_l326_c3_97ed_cond : unsigned(0 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_97ed_iftrue : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_97ed_iffalse : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_97ed_return_output : unsigned(7 downto 0);

-- layer0_node29_MUX[bit_math_h_l337_c3_7a23]
signal layer0_node29_MUX_bit_math_h_l337_c3_7a23_cond : unsigned(0 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_7a23_iftrue : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_7a23_iffalse : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_7a23_return_output : unsigned(7 downto 0);

-- layer0_node30_MUX[bit_math_h_l348_c3_7ed3]
signal layer0_node30_MUX_bit_math_h_l348_c3_7ed3_cond : unsigned(0 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iftrue : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iffalse : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_7ed3_return_output : unsigned(7 downto 0);

-- layer0_node31_MUX[bit_math_h_l359_c3_208c]
signal layer0_node31_MUX_bit_math_h_l359_c3_208c_cond : unsigned(0 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_208c_iftrue : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_208c_iffalse : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_208c_return_output : unsigned(7 downto 0);

-- layer0_node32_MUX[bit_math_h_l370_c3_bcd8]
signal layer0_node32_MUX_bit_math_h_l370_c3_bcd8_cond : unsigned(0 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iftrue : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iffalse : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_bcd8_return_output : unsigned(7 downto 0);

-- layer0_node33_MUX[bit_math_h_l381_c3_0aac]
signal layer0_node33_MUX_bit_math_h_l381_c3_0aac_cond : unsigned(0 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_0aac_iftrue : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_0aac_iffalse : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_0aac_return_output : unsigned(7 downto 0);

-- layer0_node34_MUX[bit_math_h_l392_c3_6801]
signal layer0_node34_MUX_bit_math_h_l392_c3_6801_cond : unsigned(0 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_6801_iftrue : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_6801_iffalse : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_6801_return_output : unsigned(7 downto 0);

-- layer0_node35_MUX[bit_math_h_l403_c3_749b]
signal layer0_node35_MUX_bit_math_h_l403_c3_749b_cond : unsigned(0 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_749b_iftrue : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_749b_iffalse : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_749b_return_output : unsigned(7 downto 0);

-- layer0_node36_MUX[bit_math_h_l414_c3_0db7]
signal layer0_node36_MUX_bit_math_h_l414_c3_0db7_cond : unsigned(0 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_0db7_iftrue : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_0db7_iffalse : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_0db7_return_output : unsigned(7 downto 0);

-- layer0_node37_MUX[bit_math_h_l425_c3_7f65]
signal layer0_node37_MUX_bit_math_h_l425_c3_7f65_cond : unsigned(0 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_7f65_iftrue : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_7f65_iffalse : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_7f65_return_output : unsigned(7 downto 0);

-- layer0_node38_MUX[bit_math_h_l436_c3_d774]
signal layer0_node38_MUX_bit_math_h_l436_c3_d774_cond : unsigned(0 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_d774_iftrue : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_d774_iffalse : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_d774_return_output : unsigned(7 downto 0);

-- layer0_node39_MUX[bit_math_h_l447_c3_b0c4]
signal layer0_node39_MUX_bit_math_h_l447_c3_b0c4_cond : unsigned(0 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iftrue : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iffalse : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_b0c4_return_output : unsigned(7 downto 0);

-- layer0_node40_MUX[bit_math_h_l458_c3_773e]
signal layer0_node40_MUX_bit_math_h_l458_c3_773e_cond : unsigned(0 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_773e_iftrue : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_773e_iffalse : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_773e_return_output : unsigned(7 downto 0);

-- layer0_node41_MUX[bit_math_h_l469_c3_62cc]
signal layer0_node41_MUX_bit_math_h_l469_c3_62cc_cond : unsigned(0 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_62cc_iftrue : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_62cc_iffalse : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_62cc_return_output : unsigned(7 downto 0);

-- layer0_node42_MUX[bit_math_h_l480_c3_d626]
signal layer0_node42_MUX_bit_math_h_l480_c3_d626_cond : unsigned(0 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_d626_iftrue : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_d626_iffalse : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_d626_return_output : unsigned(7 downto 0);

-- layer0_node43_MUX[bit_math_h_l491_c3_001b]
signal layer0_node43_MUX_bit_math_h_l491_c3_001b_cond : unsigned(0 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_001b_iftrue : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_001b_iffalse : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_001b_return_output : unsigned(7 downto 0);

-- layer0_node44_MUX[bit_math_h_l502_c3_1816]
signal layer0_node44_MUX_bit_math_h_l502_c3_1816_cond : unsigned(0 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_1816_iftrue : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_1816_iffalse : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_1816_return_output : unsigned(7 downto 0);

-- layer0_node45_MUX[bit_math_h_l513_c3_cc83]
signal layer0_node45_MUX_bit_math_h_l513_c3_cc83_cond : unsigned(0 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_cc83_iftrue : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_cc83_iffalse : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_cc83_return_output : unsigned(7 downto 0);

-- layer0_node46_MUX[bit_math_h_l524_c3_aa0a]
signal layer0_node46_MUX_bit_math_h_l524_c3_aa0a_cond : unsigned(0 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iftrue : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iffalse : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_aa0a_return_output : unsigned(7 downto 0);

-- layer0_node47_MUX[bit_math_h_l535_c3_167a]
signal layer0_node47_MUX_bit_math_h_l535_c3_167a_cond : unsigned(0 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_167a_iftrue : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_167a_iffalse : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_167a_return_output : unsigned(7 downto 0);

-- layer0_node48_MUX[bit_math_h_l546_c3_41a2]
signal layer0_node48_MUX_bit_math_h_l546_c3_41a2_cond : unsigned(0 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_41a2_iftrue : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_41a2_iffalse : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_41a2_return_output : unsigned(7 downto 0);

-- layer0_node49_MUX[bit_math_h_l557_c3_3c6d]
signal layer0_node49_MUX_bit_math_h_l557_c3_3c6d_cond : unsigned(0 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iftrue : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iffalse : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_3c6d_return_output : unsigned(7 downto 0);

-- layer0_node50_MUX[bit_math_h_l568_c3_e0e2]
signal layer0_node50_MUX_bit_math_h_l568_c3_e0e2_cond : unsigned(0 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iftrue : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iffalse : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_e0e2_return_output : unsigned(7 downto 0);

-- layer0_node51_MUX[bit_math_h_l579_c3_1b2f]
signal layer0_node51_MUX_bit_math_h_l579_c3_1b2f_cond : unsigned(0 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iftrue : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iffalse : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_1b2f_return_output : unsigned(7 downto 0);

-- layer0_node52_MUX[bit_math_h_l590_c3_dee1]
signal layer0_node52_MUX_bit_math_h_l590_c3_dee1_cond : unsigned(0 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_dee1_iftrue : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_dee1_iffalse : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_dee1_return_output : unsigned(7 downto 0);

-- layer0_node53_MUX[bit_math_h_l601_c3_76ac]
signal layer0_node53_MUX_bit_math_h_l601_c3_76ac_cond : unsigned(0 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_76ac_iftrue : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_76ac_iffalse : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_76ac_return_output : unsigned(7 downto 0);

-- layer0_node54_MUX[bit_math_h_l612_c3_e1c8]
signal layer0_node54_MUX_bit_math_h_l612_c3_e1c8_cond : unsigned(0 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iftrue : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iffalse : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_e1c8_return_output : unsigned(7 downto 0);

-- layer0_node55_MUX[bit_math_h_l623_c3_ec7e]
signal layer0_node55_MUX_bit_math_h_l623_c3_ec7e_cond : unsigned(0 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iftrue : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iffalse : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_ec7e_return_output : unsigned(7 downto 0);

-- layer0_node56_MUX[bit_math_h_l634_c3_5b10]
signal layer0_node56_MUX_bit_math_h_l634_c3_5b10_cond : unsigned(0 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_5b10_iftrue : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_5b10_iffalse : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_5b10_return_output : unsigned(7 downto 0);

-- layer0_node57_MUX[bit_math_h_l645_c3_d7f5]
signal layer0_node57_MUX_bit_math_h_l645_c3_d7f5_cond : unsigned(0 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iftrue : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iffalse : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_d7f5_return_output : unsigned(7 downto 0);

-- layer0_node58_MUX[bit_math_h_l656_c3_e8c0]
signal layer0_node58_MUX_bit_math_h_l656_c3_e8c0_cond : unsigned(0 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iftrue : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iffalse : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_e8c0_return_output : unsigned(7 downto 0);

-- layer0_node59_MUX[bit_math_h_l667_c3_1ea2]
signal layer0_node59_MUX_bit_math_h_l667_c3_1ea2_cond : unsigned(0 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iftrue : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iffalse : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_1ea2_return_output : unsigned(7 downto 0);

-- layer0_node60_MUX[bit_math_h_l678_c3_fe9f]
signal layer0_node60_MUX_bit_math_h_l678_c3_fe9f_cond : unsigned(0 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iftrue : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iffalse : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_fe9f_return_output : unsigned(7 downto 0);

-- layer0_node61_MUX[bit_math_h_l689_c3_9f98]
signal layer0_node61_MUX_bit_math_h_l689_c3_9f98_cond : unsigned(0 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_9f98_iftrue : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_9f98_iffalse : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_9f98_return_output : unsigned(7 downto 0);

-- layer0_node62_MUX[bit_math_h_l700_c3_0d13]
signal layer0_node62_MUX_bit_math_h_l700_c3_0d13_cond : unsigned(0 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_0d13_iftrue : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_0d13_iffalse : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_0d13_return_output : unsigned(7 downto 0);

-- layer0_node63_MUX[bit_math_h_l711_c3_2778]
signal layer0_node63_MUX_bit_math_h_l711_c3_2778_cond : unsigned(0 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_2778_iftrue : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_2778_iffalse : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_2778_return_output : unsigned(7 downto 0);

-- layer1_node0_MUX[bit_math_h_l728_c3_67cd]
signal layer1_node0_MUX_bit_math_h_l728_c3_67cd_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_67cd_iftrue : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_67cd_iffalse : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_67cd_return_output : unsigned(7 downto 0);

-- layer1_node1_MUX[bit_math_h_l739_c3_5e54]
signal layer1_node1_MUX_bit_math_h_l739_c3_5e54_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_5e54_iftrue : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_5e54_iffalse : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_5e54_return_output : unsigned(7 downto 0);

-- layer1_node2_MUX[bit_math_h_l750_c3_386d]
signal layer1_node2_MUX_bit_math_h_l750_c3_386d_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_386d_iftrue : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_386d_iffalse : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_386d_return_output : unsigned(7 downto 0);

-- layer1_node3_MUX[bit_math_h_l761_c3_c96d]
signal layer1_node3_MUX_bit_math_h_l761_c3_c96d_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_c96d_iftrue : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_c96d_iffalse : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_c96d_return_output : unsigned(7 downto 0);

-- layer1_node4_MUX[bit_math_h_l772_c3_535b]
signal layer1_node4_MUX_bit_math_h_l772_c3_535b_cond : unsigned(0 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_535b_iftrue : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_535b_iffalse : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_535b_return_output : unsigned(7 downto 0);

-- layer1_node5_MUX[bit_math_h_l783_c3_7132]
signal layer1_node5_MUX_bit_math_h_l783_c3_7132_cond : unsigned(0 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_7132_iftrue : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_7132_iffalse : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_7132_return_output : unsigned(7 downto 0);

-- layer1_node6_MUX[bit_math_h_l794_c3_59a7]
signal layer1_node6_MUX_bit_math_h_l794_c3_59a7_cond : unsigned(0 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_59a7_iftrue : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_59a7_iffalse : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_59a7_return_output : unsigned(7 downto 0);

-- layer1_node7_MUX[bit_math_h_l805_c3_a7b7]
signal layer1_node7_MUX_bit_math_h_l805_c3_a7b7_cond : unsigned(0 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iftrue : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iffalse : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_a7b7_return_output : unsigned(7 downto 0);

-- layer1_node8_MUX[bit_math_h_l816_c3_7279]
signal layer1_node8_MUX_bit_math_h_l816_c3_7279_cond : unsigned(0 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_7279_iftrue : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_7279_iffalse : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_7279_return_output : unsigned(7 downto 0);

-- layer1_node9_MUX[bit_math_h_l827_c3_90fc]
signal layer1_node9_MUX_bit_math_h_l827_c3_90fc_cond : unsigned(0 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_90fc_iftrue : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_90fc_iffalse : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_90fc_return_output : unsigned(7 downto 0);

-- layer1_node10_MUX[bit_math_h_l838_c3_e624]
signal layer1_node10_MUX_bit_math_h_l838_c3_e624_cond : unsigned(0 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_e624_iftrue : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_e624_iffalse : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_e624_return_output : unsigned(7 downto 0);

-- layer1_node11_MUX[bit_math_h_l849_c3_0669]
signal layer1_node11_MUX_bit_math_h_l849_c3_0669_cond : unsigned(0 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_0669_iftrue : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_0669_iffalse : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_0669_return_output : unsigned(7 downto 0);

-- layer1_node12_MUX[bit_math_h_l860_c3_f017]
signal layer1_node12_MUX_bit_math_h_l860_c3_f017_cond : unsigned(0 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_f017_iftrue : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_f017_iffalse : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_f017_return_output : unsigned(7 downto 0);

-- layer1_node13_MUX[bit_math_h_l871_c3_9f0e]
signal layer1_node13_MUX_bit_math_h_l871_c3_9f0e_cond : unsigned(0 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iftrue : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iffalse : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_9f0e_return_output : unsigned(7 downto 0);

-- layer1_node14_MUX[bit_math_h_l882_c3_9be0]
signal layer1_node14_MUX_bit_math_h_l882_c3_9be0_cond : unsigned(0 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_9be0_iftrue : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_9be0_iffalse : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_9be0_return_output : unsigned(7 downto 0);

-- layer1_node15_MUX[bit_math_h_l893_c3_db88]
signal layer1_node15_MUX_bit_math_h_l893_c3_db88_cond : unsigned(0 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_db88_iftrue : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_db88_iffalse : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_db88_return_output : unsigned(7 downto 0);

-- layer1_node16_MUX[bit_math_h_l904_c3_fdb3]
signal layer1_node16_MUX_bit_math_h_l904_c3_fdb3_cond : unsigned(0 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iftrue : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iffalse : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_fdb3_return_output : unsigned(7 downto 0);

-- layer1_node17_MUX[bit_math_h_l915_c3_bba5]
signal layer1_node17_MUX_bit_math_h_l915_c3_bba5_cond : unsigned(0 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_bba5_iftrue : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_bba5_iffalse : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_bba5_return_output : unsigned(7 downto 0);

-- layer1_node18_MUX[bit_math_h_l926_c3_ab1a]
signal layer1_node18_MUX_bit_math_h_l926_c3_ab1a_cond : unsigned(0 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iftrue : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iffalse : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_ab1a_return_output : unsigned(7 downto 0);

-- layer1_node19_MUX[bit_math_h_l937_c3_1a24]
signal layer1_node19_MUX_bit_math_h_l937_c3_1a24_cond : unsigned(0 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_1a24_iftrue : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_1a24_iffalse : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_1a24_return_output : unsigned(7 downto 0);

-- layer1_node20_MUX[bit_math_h_l948_c3_2dbc]
signal layer1_node20_MUX_bit_math_h_l948_c3_2dbc_cond : unsigned(0 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iftrue : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iffalse : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2dbc_return_output : unsigned(7 downto 0);

-- layer1_node21_MUX[bit_math_h_l959_c3_f718]
signal layer1_node21_MUX_bit_math_h_l959_c3_f718_cond : unsigned(0 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_f718_iftrue : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_f718_iffalse : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_f718_return_output : unsigned(7 downto 0);

-- layer1_node22_MUX[bit_math_h_l970_c3_3aa5]
signal layer1_node22_MUX_bit_math_h_l970_c3_3aa5_cond : unsigned(0 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iftrue : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iffalse : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_3aa5_return_output : unsigned(7 downto 0);

-- layer1_node23_MUX[bit_math_h_l981_c3_d2b9]
signal layer1_node23_MUX_bit_math_h_l981_c3_d2b9_cond : unsigned(0 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iftrue : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iffalse : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_d2b9_return_output : unsigned(7 downto 0);

-- layer1_node24_MUX[bit_math_h_l992_c3_8792]
signal layer1_node24_MUX_bit_math_h_l992_c3_8792_cond : unsigned(0 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_8792_iftrue : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_8792_iffalse : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_8792_return_output : unsigned(7 downto 0);

-- layer1_node25_MUX[bit_math_h_l1003_c3_2c90]
signal layer1_node25_MUX_bit_math_h_l1003_c3_2c90_cond : unsigned(0 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iftrue : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iffalse : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_2c90_return_output : unsigned(7 downto 0);

-- layer1_node26_MUX[bit_math_h_l1014_c3_f8c1]
signal layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_cond : unsigned(0 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iftrue : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iffalse : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_return_output : unsigned(7 downto 0);

-- layer1_node27_MUX[bit_math_h_l1025_c3_7ac4]
signal layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_cond : unsigned(0 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iftrue : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iffalse : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_return_output : unsigned(7 downto 0);

-- layer1_node28_MUX[bit_math_h_l1036_c3_deef]
signal layer1_node28_MUX_bit_math_h_l1036_c3_deef_cond : unsigned(0 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_deef_iftrue : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_deef_iffalse : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_deef_return_output : unsigned(7 downto 0);

-- layer1_node29_MUX[bit_math_h_l1047_c3_d4d6]
signal layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_cond : unsigned(0 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iftrue : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iffalse : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_return_output : unsigned(7 downto 0);

-- layer1_node30_MUX[bit_math_h_l1058_c3_d1f5]
signal layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_cond : unsigned(0 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iftrue : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iffalse : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_return_output : unsigned(7 downto 0);

-- layer1_node31_MUX[bit_math_h_l1069_c3_fc71]
signal layer1_node31_MUX_bit_math_h_l1069_c3_fc71_cond : unsigned(0 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iftrue : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iffalse : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_fc71_return_output : unsigned(7 downto 0);

-- layer2_node0_MUX[bit_math_h_l1086_c3_5a52]
signal layer2_node0_MUX_bit_math_h_l1086_c3_5a52_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iftrue : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iffalse : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_5a52_return_output : unsigned(7 downto 0);

-- layer2_node1_MUX[bit_math_h_l1097_c3_fc1c]
signal layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iftrue : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iffalse : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_return_output : unsigned(7 downto 0);

-- layer2_node2_MUX[bit_math_h_l1108_c3_922a]
signal layer2_node2_MUX_bit_math_h_l1108_c3_922a_cond : unsigned(0 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_922a_iftrue : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_922a_iffalse : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_922a_return_output : unsigned(7 downto 0);

-- layer2_node3_MUX[bit_math_h_l1119_c3_b25e]
signal layer2_node3_MUX_bit_math_h_l1119_c3_b25e_cond : unsigned(0 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iftrue : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iffalse : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_b25e_return_output : unsigned(7 downto 0);

-- layer2_node4_MUX[bit_math_h_l1130_c3_5fd5]
signal layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_cond : unsigned(0 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iftrue : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iffalse : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_return_output : unsigned(7 downto 0);

-- layer2_node5_MUX[bit_math_h_l1141_c3_6ecd]
signal layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_cond : unsigned(0 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iftrue : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iffalse : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_return_output : unsigned(7 downto 0);

-- layer2_node6_MUX[bit_math_h_l1152_c3_d917]
signal layer2_node6_MUX_bit_math_h_l1152_c3_d917_cond : unsigned(0 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_d917_iftrue : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_d917_iffalse : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_d917_return_output : unsigned(7 downto 0);

-- layer2_node7_MUX[bit_math_h_l1163_c3_d44d]
signal layer2_node7_MUX_bit_math_h_l1163_c3_d44d_cond : unsigned(0 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iftrue : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iffalse : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_d44d_return_output : unsigned(7 downto 0);

-- layer2_node8_MUX[bit_math_h_l1174_c3_d504]
signal layer2_node8_MUX_bit_math_h_l1174_c3_d504_cond : unsigned(0 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_d504_iftrue : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_d504_iffalse : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_d504_return_output : unsigned(7 downto 0);

-- layer2_node9_MUX[bit_math_h_l1185_c3_8a90]
signal layer2_node9_MUX_bit_math_h_l1185_c3_8a90_cond : unsigned(0 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iftrue : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iffalse : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_8a90_return_output : unsigned(7 downto 0);

-- layer2_node10_MUX[bit_math_h_l1196_c3_c6ad]
signal layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_cond : unsigned(0 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iftrue : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iffalse : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_return_output : unsigned(7 downto 0);

-- layer2_node11_MUX[bit_math_h_l1207_c3_e593]
signal layer2_node11_MUX_bit_math_h_l1207_c3_e593_cond : unsigned(0 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_e593_iftrue : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_e593_iffalse : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_e593_return_output : unsigned(7 downto 0);

-- layer2_node12_MUX[bit_math_h_l1218_c3_ed0c]
signal layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_cond : unsigned(0 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iftrue : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iffalse : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_return_output : unsigned(7 downto 0);

-- layer2_node13_MUX[bit_math_h_l1229_c3_d88d]
signal layer2_node13_MUX_bit_math_h_l1229_c3_d88d_cond : unsigned(0 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iftrue : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iffalse : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_d88d_return_output : unsigned(7 downto 0);

-- layer2_node14_MUX[bit_math_h_l1240_c3_d3d6]
signal layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_cond : unsigned(0 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iftrue : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iffalse : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_return_output : unsigned(7 downto 0);

-- layer2_node15_MUX[bit_math_h_l1251_c3_03ac]
signal layer2_node15_MUX_bit_math_h_l1251_c3_03ac_cond : unsigned(0 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iftrue : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iffalse : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_03ac_return_output : unsigned(7 downto 0);

-- layer3_node0_MUX[bit_math_h_l1268_c3_6917]
signal layer3_node0_MUX_bit_math_h_l1268_c3_6917_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_6917_iftrue : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_6917_iffalse : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_6917_return_output : unsigned(7 downto 0);

-- layer3_node1_MUX[bit_math_h_l1279_c3_e270]
signal layer3_node1_MUX_bit_math_h_l1279_c3_e270_cond : unsigned(0 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_e270_iftrue : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_e270_iffalse : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_e270_return_output : unsigned(7 downto 0);

-- layer3_node2_MUX[bit_math_h_l1290_c3_769c]
signal layer3_node2_MUX_bit_math_h_l1290_c3_769c_cond : unsigned(0 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_769c_iftrue : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_769c_iffalse : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_769c_return_output : unsigned(7 downto 0);

-- layer3_node3_MUX[bit_math_h_l1301_c3_fb21]
signal layer3_node3_MUX_bit_math_h_l1301_c3_fb21_cond : unsigned(0 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iftrue : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iffalse : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_fb21_return_output : unsigned(7 downto 0);

-- layer3_node4_MUX[bit_math_h_l1312_c3_f274]
signal layer3_node4_MUX_bit_math_h_l1312_c3_f274_cond : unsigned(0 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_f274_iftrue : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_f274_iffalse : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_f274_return_output : unsigned(7 downto 0);

-- layer3_node5_MUX[bit_math_h_l1323_c3_6b46]
signal layer3_node5_MUX_bit_math_h_l1323_c3_6b46_cond : unsigned(0 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iftrue : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iffalse : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_6b46_return_output : unsigned(7 downto 0);

-- layer3_node6_MUX[bit_math_h_l1334_c3_41a0]
signal layer3_node6_MUX_bit_math_h_l1334_c3_41a0_cond : unsigned(0 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iftrue : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iffalse : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_41a0_return_output : unsigned(7 downto 0);

-- layer3_node7_MUX[bit_math_h_l1345_c3_969c]
signal layer3_node7_MUX_bit_math_h_l1345_c3_969c_cond : unsigned(0 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_969c_iftrue : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_969c_iffalse : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_969c_return_output : unsigned(7 downto 0);

-- layer4_node0_MUX[bit_math_h_l1362_c3_b41d]
signal layer4_node0_MUX_bit_math_h_l1362_c3_b41d_cond : unsigned(0 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iftrue : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iffalse : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_b41d_return_output : unsigned(7 downto 0);

-- layer4_node1_MUX[bit_math_h_l1373_c3_f2a6]
signal layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_cond : unsigned(0 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iftrue : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iffalse : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_return_output : unsigned(7 downto 0);

-- layer4_node2_MUX[bit_math_h_l1384_c3_3339]
signal layer4_node2_MUX_bit_math_h_l1384_c3_3339_cond : unsigned(0 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_3339_iftrue : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_3339_iffalse : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_3339_return_output : unsigned(7 downto 0);

-- layer4_node3_MUX[bit_math_h_l1395_c3_b75d]
signal layer4_node3_MUX_bit_math_h_l1395_c3_b75d_cond : unsigned(0 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iftrue : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iffalse : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_b75d_return_output : unsigned(7 downto 0);

-- layer5_node0_MUX[bit_math_h_l1412_c3_5f1f]
signal layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_cond : unsigned(0 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iftrue : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iffalse : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_return_output : unsigned(7 downto 0);

-- layer5_node1_MUX[bit_math_h_l1423_c3_1d22]
signal layer5_node1_MUX_bit_math_h_l1423_c3_1d22_cond : unsigned(0 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iftrue : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iffalse : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_1d22_return_output : unsigned(7 downto 0);

-- layer6_node0_MUX[bit_math_h_l1440_c3_247e]
signal layer6_node0_MUX_bit_math_h_l1440_c3_247e_cond : unsigned(0 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_247e_iftrue : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_247e_iffalse : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_247e_return_output : unsigned(7 downto 0);

function uint7_0_0( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint7_1_1( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint7_2_2( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint7_3_3( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;

function uint7_4_4( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(4- i);
      end loop;
return return_output;
end function;

function uint7_5_5( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(5- i);
      end loop;
return return_output;
end function;

function uint7_6_6( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(6- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_8bd4
layer0_node0_MUX_bit_math_h_l18_c3_8bd4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_8bd4_cond,
layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_8bd4_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_b2fc
layer0_node1_MUX_bit_math_h_l29_c3_b2fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_b2fc_cond,
layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_b2fc_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_3d12
layer0_node2_MUX_bit_math_h_l40_c3_3d12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_3d12_cond,
layer0_node2_MUX_bit_math_h_l40_c3_3d12_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_3d12_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_3d12_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_13b9
layer0_node3_MUX_bit_math_h_l51_c3_13b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_13b9_cond,
layer0_node3_MUX_bit_math_h_l51_c3_13b9_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_13b9_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_13b9_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_be4c
layer0_node4_MUX_bit_math_h_l62_c3_be4c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_be4c_cond,
layer0_node4_MUX_bit_math_h_l62_c3_be4c_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_be4c_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_be4c_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_936b
layer0_node5_MUX_bit_math_h_l73_c3_936b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_936b_cond,
layer0_node5_MUX_bit_math_h_l73_c3_936b_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_936b_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_936b_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_6f9a
layer0_node6_MUX_bit_math_h_l84_c3_6f9a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_6f9a_cond,
layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_6f9a_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_f259
layer0_node7_MUX_bit_math_h_l95_c3_f259 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_f259_cond,
layer0_node7_MUX_bit_math_h_l95_c3_f259_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_f259_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_f259_return_output);

-- layer0_node8_MUX_bit_math_h_l106_c3_2e0c
layer0_node8_MUX_bit_math_h_l106_c3_2e0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node8_MUX_bit_math_h_l106_c3_2e0c_cond,
layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iftrue,
layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iffalse,
layer0_node8_MUX_bit_math_h_l106_c3_2e0c_return_output);

-- layer0_node9_MUX_bit_math_h_l117_c3_1a47
layer0_node9_MUX_bit_math_h_l117_c3_1a47 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node9_MUX_bit_math_h_l117_c3_1a47_cond,
layer0_node9_MUX_bit_math_h_l117_c3_1a47_iftrue,
layer0_node9_MUX_bit_math_h_l117_c3_1a47_iffalse,
layer0_node9_MUX_bit_math_h_l117_c3_1a47_return_output);

-- layer0_node10_MUX_bit_math_h_l128_c3_0e40
layer0_node10_MUX_bit_math_h_l128_c3_0e40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node10_MUX_bit_math_h_l128_c3_0e40_cond,
layer0_node10_MUX_bit_math_h_l128_c3_0e40_iftrue,
layer0_node10_MUX_bit_math_h_l128_c3_0e40_iffalse,
layer0_node10_MUX_bit_math_h_l128_c3_0e40_return_output);

-- layer0_node11_MUX_bit_math_h_l139_c3_381c
layer0_node11_MUX_bit_math_h_l139_c3_381c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node11_MUX_bit_math_h_l139_c3_381c_cond,
layer0_node11_MUX_bit_math_h_l139_c3_381c_iftrue,
layer0_node11_MUX_bit_math_h_l139_c3_381c_iffalse,
layer0_node11_MUX_bit_math_h_l139_c3_381c_return_output);

-- layer0_node12_MUX_bit_math_h_l150_c3_1560
layer0_node12_MUX_bit_math_h_l150_c3_1560 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node12_MUX_bit_math_h_l150_c3_1560_cond,
layer0_node12_MUX_bit_math_h_l150_c3_1560_iftrue,
layer0_node12_MUX_bit_math_h_l150_c3_1560_iffalse,
layer0_node12_MUX_bit_math_h_l150_c3_1560_return_output);

-- layer0_node13_MUX_bit_math_h_l161_c3_3a1c
layer0_node13_MUX_bit_math_h_l161_c3_3a1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node13_MUX_bit_math_h_l161_c3_3a1c_cond,
layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iftrue,
layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iffalse,
layer0_node13_MUX_bit_math_h_l161_c3_3a1c_return_output);

-- layer0_node14_MUX_bit_math_h_l172_c3_7ef7
layer0_node14_MUX_bit_math_h_l172_c3_7ef7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node14_MUX_bit_math_h_l172_c3_7ef7_cond,
layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iftrue,
layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iffalse,
layer0_node14_MUX_bit_math_h_l172_c3_7ef7_return_output);

-- layer0_node15_MUX_bit_math_h_l183_c3_392b
layer0_node15_MUX_bit_math_h_l183_c3_392b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node15_MUX_bit_math_h_l183_c3_392b_cond,
layer0_node15_MUX_bit_math_h_l183_c3_392b_iftrue,
layer0_node15_MUX_bit_math_h_l183_c3_392b_iffalse,
layer0_node15_MUX_bit_math_h_l183_c3_392b_return_output);

-- layer0_node16_MUX_bit_math_h_l194_c3_cada
layer0_node16_MUX_bit_math_h_l194_c3_cada : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node16_MUX_bit_math_h_l194_c3_cada_cond,
layer0_node16_MUX_bit_math_h_l194_c3_cada_iftrue,
layer0_node16_MUX_bit_math_h_l194_c3_cada_iffalse,
layer0_node16_MUX_bit_math_h_l194_c3_cada_return_output);

-- layer0_node17_MUX_bit_math_h_l205_c3_39fd
layer0_node17_MUX_bit_math_h_l205_c3_39fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node17_MUX_bit_math_h_l205_c3_39fd_cond,
layer0_node17_MUX_bit_math_h_l205_c3_39fd_iftrue,
layer0_node17_MUX_bit_math_h_l205_c3_39fd_iffalse,
layer0_node17_MUX_bit_math_h_l205_c3_39fd_return_output);

-- layer0_node18_MUX_bit_math_h_l216_c3_23c8
layer0_node18_MUX_bit_math_h_l216_c3_23c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node18_MUX_bit_math_h_l216_c3_23c8_cond,
layer0_node18_MUX_bit_math_h_l216_c3_23c8_iftrue,
layer0_node18_MUX_bit_math_h_l216_c3_23c8_iffalse,
layer0_node18_MUX_bit_math_h_l216_c3_23c8_return_output);

-- layer0_node19_MUX_bit_math_h_l227_c3_ea58
layer0_node19_MUX_bit_math_h_l227_c3_ea58 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node19_MUX_bit_math_h_l227_c3_ea58_cond,
layer0_node19_MUX_bit_math_h_l227_c3_ea58_iftrue,
layer0_node19_MUX_bit_math_h_l227_c3_ea58_iffalse,
layer0_node19_MUX_bit_math_h_l227_c3_ea58_return_output);

-- layer0_node20_MUX_bit_math_h_l238_c3_eb78
layer0_node20_MUX_bit_math_h_l238_c3_eb78 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node20_MUX_bit_math_h_l238_c3_eb78_cond,
layer0_node20_MUX_bit_math_h_l238_c3_eb78_iftrue,
layer0_node20_MUX_bit_math_h_l238_c3_eb78_iffalse,
layer0_node20_MUX_bit_math_h_l238_c3_eb78_return_output);

-- layer0_node21_MUX_bit_math_h_l249_c3_228d
layer0_node21_MUX_bit_math_h_l249_c3_228d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node21_MUX_bit_math_h_l249_c3_228d_cond,
layer0_node21_MUX_bit_math_h_l249_c3_228d_iftrue,
layer0_node21_MUX_bit_math_h_l249_c3_228d_iffalse,
layer0_node21_MUX_bit_math_h_l249_c3_228d_return_output);

-- layer0_node22_MUX_bit_math_h_l260_c3_1c3c
layer0_node22_MUX_bit_math_h_l260_c3_1c3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node22_MUX_bit_math_h_l260_c3_1c3c_cond,
layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iftrue,
layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iffalse,
layer0_node22_MUX_bit_math_h_l260_c3_1c3c_return_output);

-- layer0_node23_MUX_bit_math_h_l271_c3_6340
layer0_node23_MUX_bit_math_h_l271_c3_6340 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node23_MUX_bit_math_h_l271_c3_6340_cond,
layer0_node23_MUX_bit_math_h_l271_c3_6340_iftrue,
layer0_node23_MUX_bit_math_h_l271_c3_6340_iffalse,
layer0_node23_MUX_bit_math_h_l271_c3_6340_return_output);

-- layer0_node24_MUX_bit_math_h_l282_c3_670b
layer0_node24_MUX_bit_math_h_l282_c3_670b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node24_MUX_bit_math_h_l282_c3_670b_cond,
layer0_node24_MUX_bit_math_h_l282_c3_670b_iftrue,
layer0_node24_MUX_bit_math_h_l282_c3_670b_iffalse,
layer0_node24_MUX_bit_math_h_l282_c3_670b_return_output);

-- layer0_node25_MUX_bit_math_h_l293_c3_83e8
layer0_node25_MUX_bit_math_h_l293_c3_83e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node25_MUX_bit_math_h_l293_c3_83e8_cond,
layer0_node25_MUX_bit_math_h_l293_c3_83e8_iftrue,
layer0_node25_MUX_bit_math_h_l293_c3_83e8_iffalse,
layer0_node25_MUX_bit_math_h_l293_c3_83e8_return_output);

-- layer0_node26_MUX_bit_math_h_l304_c3_53e2
layer0_node26_MUX_bit_math_h_l304_c3_53e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node26_MUX_bit_math_h_l304_c3_53e2_cond,
layer0_node26_MUX_bit_math_h_l304_c3_53e2_iftrue,
layer0_node26_MUX_bit_math_h_l304_c3_53e2_iffalse,
layer0_node26_MUX_bit_math_h_l304_c3_53e2_return_output);

-- layer0_node27_MUX_bit_math_h_l315_c3_ac24
layer0_node27_MUX_bit_math_h_l315_c3_ac24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node27_MUX_bit_math_h_l315_c3_ac24_cond,
layer0_node27_MUX_bit_math_h_l315_c3_ac24_iftrue,
layer0_node27_MUX_bit_math_h_l315_c3_ac24_iffalse,
layer0_node27_MUX_bit_math_h_l315_c3_ac24_return_output);

-- layer0_node28_MUX_bit_math_h_l326_c3_97ed
layer0_node28_MUX_bit_math_h_l326_c3_97ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node28_MUX_bit_math_h_l326_c3_97ed_cond,
layer0_node28_MUX_bit_math_h_l326_c3_97ed_iftrue,
layer0_node28_MUX_bit_math_h_l326_c3_97ed_iffalse,
layer0_node28_MUX_bit_math_h_l326_c3_97ed_return_output);

-- layer0_node29_MUX_bit_math_h_l337_c3_7a23
layer0_node29_MUX_bit_math_h_l337_c3_7a23 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node29_MUX_bit_math_h_l337_c3_7a23_cond,
layer0_node29_MUX_bit_math_h_l337_c3_7a23_iftrue,
layer0_node29_MUX_bit_math_h_l337_c3_7a23_iffalse,
layer0_node29_MUX_bit_math_h_l337_c3_7a23_return_output);

-- layer0_node30_MUX_bit_math_h_l348_c3_7ed3
layer0_node30_MUX_bit_math_h_l348_c3_7ed3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node30_MUX_bit_math_h_l348_c3_7ed3_cond,
layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iftrue,
layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iffalse,
layer0_node30_MUX_bit_math_h_l348_c3_7ed3_return_output);

-- layer0_node31_MUX_bit_math_h_l359_c3_208c
layer0_node31_MUX_bit_math_h_l359_c3_208c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node31_MUX_bit_math_h_l359_c3_208c_cond,
layer0_node31_MUX_bit_math_h_l359_c3_208c_iftrue,
layer0_node31_MUX_bit_math_h_l359_c3_208c_iffalse,
layer0_node31_MUX_bit_math_h_l359_c3_208c_return_output);

-- layer0_node32_MUX_bit_math_h_l370_c3_bcd8
layer0_node32_MUX_bit_math_h_l370_c3_bcd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node32_MUX_bit_math_h_l370_c3_bcd8_cond,
layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iftrue,
layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iffalse,
layer0_node32_MUX_bit_math_h_l370_c3_bcd8_return_output);

-- layer0_node33_MUX_bit_math_h_l381_c3_0aac
layer0_node33_MUX_bit_math_h_l381_c3_0aac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node33_MUX_bit_math_h_l381_c3_0aac_cond,
layer0_node33_MUX_bit_math_h_l381_c3_0aac_iftrue,
layer0_node33_MUX_bit_math_h_l381_c3_0aac_iffalse,
layer0_node33_MUX_bit_math_h_l381_c3_0aac_return_output);

-- layer0_node34_MUX_bit_math_h_l392_c3_6801
layer0_node34_MUX_bit_math_h_l392_c3_6801 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node34_MUX_bit_math_h_l392_c3_6801_cond,
layer0_node34_MUX_bit_math_h_l392_c3_6801_iftrue,
layer0_node34_MUX_bit_math_h_l392_c3_6801_iffalse,
layer0_node34_MUX_bit_math_h_l392_c3_6801_return_output);

-- layer0_node35_MUX_bit_math_h_l403_c3_749b
layer0_node35_MUX_bit_math_h_l403_c3_749b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node35_MUX_bit_math_h_l403_c3_749b_cond,
layer0_node35_MUX_bit_math_h_l403_c3_749b_iftrue,
layer0_node35_MUX_bit_math_h_l403_c3_749b_iffalse,
layer0_node35_MUX_bit_math_h_l403_c3_749b_return_output);

-- layer0_node36_MUX_bit_math_h_l414_c3_0db7
layer0_node36_MUX_bit_math_h_l414_c3_0db7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node36_MUX_bit_math_h_l414_c3_0db7_cond,
layer0_node36_MUX_bit_math_h_l414_c3_0db7_iftrue,
layer0_node36_MUX_bit_math_h_l414_c3_0db7_iffalse,
layer0_node36_MUX_bit_math_h_l414_c3_0db7_return_output);

-- layer0_node37_MUX_bit_math_h_l425_c3_7f65
layer0_node37_MUX_bit_math_h_l425_c3_7f65 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node37_MUX_bit_math_h_l425_c3_7f65_cond,
layer0_node37_MUX_bit_math_h_l425_c3_7f65_iftrue,
layer0_node37_MUX_bit_math_h_l425_c3_7f65_iffalse,
layer0_node37_MUX_bit_math_h_l425_c3_7f65_return_output);

-- layer0_node38_MUX_bit_math_h_l436_c3_d774
layer0_node38_MUX_bit_math_h_l436_c3_d774 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node38_MUX_bit_math_h_l436_c3_d774_cond,
layer0_node38_MUX_bit_math_h_l436_c3_d774_iftrue,
layer0_node38_MUX_bit_math_h_l436_c3_d774_iffalse,
layer0_node38_MUX_bit_math_h_l436_c3_d774_return_output);

-- layer0_node39_MUX_bit_math_h_l447_c3_b0c4
layer0_node39_MUX_bit_math_h_l447_c3_b0c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node39_MUX_bit_math_h_l447_c3_b0c4_cond,
layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iftrue,
layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iffalse,
layer0_node39_MUX_bit_math_h_l447_c3_b0c4_return_output);

-- layer0_node40_MUX_bit_math_h_l458_c3_773e
layer0_node40_MUX_bit_math_h_l458_c3_773e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node40_MUX_bit_math_h_l458_c3_773e_cond,
layer0_node40_MUX_bit_math_h_l458_c3_773e_iftrue,
layer0_node40_MUX_bit_math_h_l458_c3_773e_iffalse,
layer0_node40_MUX_bit_math_h_l458_c3_773e_return_output);

-- layer0_node41_MUX_bit_math_h_l469_c3_62cc
layer0_node41_MUX_bit_math_h_l469_c3_62cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node41_MUX_bit_math_h_l469_c3_62cc_cond,
layer0_node41_MUX_bit_math_h_l469_c3_62cc_iftrue,
layer0_node41_MUX_bit_math_h_l469_c3_62cc_iffalse,
layer0_node41_MUX_bit_math_h_l469_c3_62cc_return_output);

-- layer0_node42_MUX_bit_math_h_l480_c3_d626
layer0_node42_MUX_bit_math_h_l480_c3_d626 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node42_MUX_bit_math_h_l480_c3_d626_cond,
layer0_node42_MUX_bit_math_h_l480_c3_d626_iftrue,
layer0_node42_MUX_bit_math_h_l480_c3_d626_iffalse,
layer0_node42_MUX_bit_math_h_l480_c3_d626_return_output);

-- layer0_node43_MUX_bit_math_h_l491_c3_001b
layer0_node43_MUX_bit_math_h_l491_c3_001b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node43_MUX_bit_math_h_l491_c3_001b_cond,
layer0_node43_MUX_bit_math_h_l491_c3_001b_iftrue,
layer0_node43_MUX_bit_math_h_l491_c3_001b_iffalse,
layer0_node43_MUX_bit_math_h_l491_c3_001b_return_output);

-- layer0_node44_MUX_bit_math_h_l502_c3_1816
layer0_node44_MUX_bit_math_h_l502_c3_1816 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node44_MUX_bit_math_h_l502_c3_1816_cond,
layer0_node44_MUX_bit_math_h_l502_c3_1816_iftrue,
layer0_node44_MUX_bit_math_h_l502_c3_1816_iffalse,
layer0_node44_MUX_bit_math_h_l502_c3_1816_return_output);

-- layer0_node45_MUX_bit_math_h_l513_c3_cc83
layer0_node45_MUX_bit_math_h_l513_c3_cc83 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node45_MUX_bit_math_h_l513_c3_cc83_cond,
layer0_node45_MUX_bit_math_h_l513_c3_cc83_iftrue,
layer0_node45_MUX_bit_math_h_l513_c3_cc83_iffalse,
layer0_node45_MUX_bit_math_h_l513_c3_cc83_return_output);

-- layer0_node46_MUX_bit_math_h_l524_c3_aa0a
layer0_node46_MUX_bit_math_h_l524_c3_aa0a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node46_MUX_bit_math_h_l524_c3_aa0a_cond,
layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iftrue,
layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iffalse,
layer0_node46_MUX_bit_math_h_l524_c3_aa0a_return_output);

-- layer0_node47_MUX_bit_math_h_l535_c3_167a
layer0_node47_MUX_bit_math_h_l535_c3_167a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node47_MUX_bit_math_h_l535_c3_167a_cond,
layer0_node47_MUX_bit_math_h_l535_c3_167a_iftrue,
layer0_node47_MUX_bit_math_h_l535_c3_167a_iffalse,
layer0_node47_MUX_bit_math_h_l535_c3_167a_return_output);

-- layer0_node48_MUX_bit_math_h_l546_c3_41a2
layer0_node48_MUX_bit_math_h_l546_c3_41a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node48_MUX_bit_math_h_l546_c3_41a2_cond,
layer0_node48_MUX_bit_math_h_l546_c3_41a2_iftrue,
layer0_node48_MUX_bit_math_h_l546_c3_41a2_iffalse,
layer0_node48_MUX_bit_math_h_l546_c3_41a2_return_output);

-- layer0_node49_MUX_bit_math_h_l557_c3_3c6d
layer0_node49_MUX_bit_math_h_l557_c3_3c6d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node49_MUX_bit_math_h_l557_c3_3c6d_cond,
layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iftrue,
layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iffalse,
layer0_node49_MUX_bit_math_h_l557_c3_3c6d_return_output);

-- layer0_node50_MUX_bit_math_h_l568_c3_e0e2
layer0_node50_MUX_bit_math_h_l568_c3_e0e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node50_MUX_bit_math_h_l568_c3_e0e2_cond,
layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iftrue,
layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iffalse,
layer0_node50_MUX_bit_math_h_l568_c3_e0e2_return_output);

-- layer0_node51_MUX_bit_math_h_l579_c3_1b2f
layer0_node51_MUX_bit_math_h_l579_c3_1b2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node51_MUX_bit_math_h_l579_c3_1b2f_cond,
layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iftrue,
layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iffalse,
layer0_node51_MUX_bit_math_h_l579_c3_1b2f_return_output);

-- layer0_node52_MUX_bit_math_h_l590_c3_dee1
layer0_node52_MUX_bit_math_h_l590_c3_dee1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node52_MUX_bit_math_h_l590_c3_dee1_cond,
layer0_node52_MUX_bit_math_h_l590_c3_dee1_iftrue,
layer0_node52_MUX_bit_math_h_l590_c3_dee1_iffalse,
layer0_node52_MUX_bit_math_h_l590_c3_dee1_return_output);

-- layer0_node53_MUX_bit_math_h_l601_c3_76ac
layer0_node53_MUX_bit_math_h_l601_c3_76ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node53_MUX_bit_math_h_l601_c3_76ac_cond,
layer0_node53_MUX_bit_math_h_l601_c3_76ac_iftrue,
layer0_node53_MUX_bit_math_h_l601_c3_76ac_iffalse,
layer0_node53_MUX_bit_math_h_l601_c3_76ac_return_output);

-- layer0_node54_MUX_bit_math_h_l612_c3_e1c8
layer0_node54_MUX_bit_math_h_l612_c3_e1c8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node54_MUX_bit_math_h_l612_c3_e1c8_cond,
layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iftrue,
layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iffalse,
layer0_node54_MUX_bit_math_h_l612_c3_e1c8_return_output);

-- layer0_node55_MUX_bit_math_h_l623_c3_ec7e
layer0_node55_MUX_bit_math_h_l623_c3_ec7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node55_MUX_bit_math_h_l623_c3_ec7e_cond,
layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iftrue,
layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iffalse,
layer0_node55_MUX_bit_math_h_l623_c3_ec7e_return_output);

-- layer0_node56_MUX_bit_math_h_l634_c3_5b10
layer0_node56_MUX_bit_math_h_l634_c3_5b10 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node56_MUX_bit_math_h_l634_c3_5b10_cond,
layer0_node56_MUX_bit_math_h_l634_c3_5b10_iftrue,
layer0_node56_MUX_bit_math_h_l634_c3_5b10_iffalse,
layer0_node56_MUX_bit_math_h_l634_c3_5b10_return_output);

-- layer0_node57_MUX_bit_math_h_l645_c3_d7f5
layer0_node57_MUX_bit_math_h_l645_c3_d7f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node57_MUX_bit_math_h_l645_c3_d7f5_cond,
layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iftrue,
layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iffalse,
layer0_node57_MUX_bit_math_h_l645_c3_d7f5_return_output);

-- layer0_node58_MUX_bit_math_h_l656_c3_e8c0
layer0_node58_MUX_bit_math_h_l656_c3_e8c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node58_MUX_bit_math_h_l656_c3_e8c0_cond,
layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iftrue,
layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iffalse,
layer0_node58_MUX_bit_math_h_l656_c3_e8c0_return_output);

-- layer0_node59_MUX_bit_math_h_l667_c3_1ea2
layer0_node59_MUX_bit_math_h_l667_c3_1ea2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node59_MUX_bit_math_h_l667_c3_1ea2_cond,
layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iftrue,
layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iffalse,
layer0_node59_MUX_bit_math_h_l667_c3_1ea2_return_output);

-- layer0_node60_MUX_bit_math_h_l678_c3_fe9f
layer0_node60_MUX_bit_math_h_l678_c3_fe9f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node60_MUX_bit_math_h_l678_c3_fe9f_cond,
layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iftrue,
layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iffalse,
layer0_node60_MUX_bit_math_h_l678_c3_fe9f_return_output);

-- layer0_node61_MUX_bit_math_h_l689_c3_9f98
layer0_node61_MUX_bit_math_h_l689_c3_9f98 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node61_MUX_bit_math_h_l689_c3_9f98_cond,
layer0_node61_MUX_bit_math_h_l689_c3_9f98_iftrue,
layer0_node61_MUX_bit_math_h_l689_c3_9f98_iffalse,
layer0_node61_MUX_bit_math_h_l689_c3_9f98_return_output);

-- layer0_node62_MUX_bit_math_h_l700_c3_0d13
layer0_node62_MUX_bit_math_h_l700_c3_0d13 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node62_MUX_bit_math_h_l700_c3_0d13_cond,
layer0_node62_MUX_bit_math_h_l700_c3_0d13_iftrue,
layer0_node62_MUX_bit_math_h_l700_c3_0d13_iffalse,
layer0_node62_MUX_bit_math_h_l700_c3_0d13_return_output);

-- layer0_node63_MUX_bit_math_h_l711_c3_2778
layer0_node63_MUX_bit_math_h_l711_c3_2778 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node63_MUX_bit_math_h_l711_c3_2778_cond,
layer0_node63_MUX_bit_math_h_l711_c3_2778_iftrue,
layer0_node63_MUX_bit_math_h_l711_c3_2778_iffalse,
layer0_node63_MUX_bit_math_h_l711_c3_2778_return_output);

-- layer1_node0_MUX_bit_math_h_l728_c3_67cd
layer1_node0_MUX_bit_math_h_l728_c3_67cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l728_c3_67cd_cond,
layer1_node0_MUX_bit_math_h_l728_c3_67cd_iftrue,
layer1_node0_MUX_bit_math_h_l728_c3_67cd_iffalse,
layer1_node0_MUX_bit_math_h_l728_c3_67cd_return_output);

-- layer1_node1_MUX_bit_math_h_l739_c3_5e54
layer1_node1_MUX_bit_math_h_l739_c3_5e54 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l739_c3_5e54_cond,
layer1_node1_MUX_bit_math_h_l739_c3_5e54_iftrue,
layer1_node1_MUX_bit_math_h_l739_c3_5e54_iffalse,
layer1_node1_MUX_bit_math_h_l739_c3_5e54_return_output);

-- layer1_node2_MUX_bit_math_h_l750_c3_386d
layer1_node2_MUX_bit_math_h_l750_c3_386d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l750_c3_386d_cond,
layer1_node2_MUX_bit_math_h_l750_c3_386d_iftrue,
layer1_node2_MUX_bit_math_h_l750_c3_386d_iffalse,
layer1_node2_MUX_bit_math_h_l750_c3_386d_return_output);

-- layer1_node3_MUX_bit_math_h_l761_c3_c96d
layer1_node3_MUX_bit_math_h_l761_c3_c96d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l761_c3_c96d_cond,
layer1_node3_MUX_bit_math_h_l761_c3_c96d_iftrue,
layer1_node3_MUX_bit_math_h_l761_c3_c96d_iffalse,
layer1_node3_MUX_bit_math_h_l761_c3_c96d_return_output);

-- layer1_node4_MUX_bit_math_h_l772_c3_535b
layer1_node4_MUX_bit_math_h_l772_c3_535b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node4_MUX_bit_math_h_l772_c3_535b_cond,
layer1_node4_MUX_bit_math_h_l772_c3_535b_iftrue,
layer1_node4_MUX_bit_math_h_l772_c3_535b_iffalse,
layer1_node4_MUX_bit_math_h_l772_c3_535b_return_output);

-- layer1_node5_MUX_bit_math_h_l783_c3_7132
layer1_node5_MUX_bit_math_h_l783_c3_7132 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node5_MUX_bit_math_h_l783_c3_7132_cond,
layer1_node5_MUX_bit_math_h_l783_c3_7132_iftrue,
layer1_node5_MUX_bit_math_h_l783_c3_7132_iffalse,
layer1_node5_MUX_bit_math_h_l783_c3_7132_return_output);

-- layer1_node6_MUX_bit_math_h_l794_c3_59a7
layer1_node6_MUX_bit_math_h_l794_c3_59a7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node6_MUX_bit_math_h_l794_c3_59a7_cond,
layer1_node6_MUX_bit_math_h_l794_c3_59a7_iftrue,
layer1_node6_MUX_bit_math_h_l794_c3_59a7_iffalse,
layer1_node6_MUX_bit_math_h_l794_c3_59a7_return_output);

-- layer1_node7_MUX_bit_math_h_l805_c3_a7b7
layer1_node7_MUX_bit_math_h_l805_c3_a7b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node7_MUX_bit_math_h_l805_c3_a7b7_cond,
layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iftrue,
layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iffalse,
layer1_node7_MUX_bit_math_h_l805_c3_a7b7_return_output);

-- layer1_node8_MUX_bit_math_h_l816_c3_7279
layer1_node8_MUX_bit_math_h_l816_c3_7279 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node8_MUX_bit_math_h_l816_c3_7279_cond,
layer1_node8_MUX_bit_math_h_l816_c3_7279_iftrue,
layer1_node8_MUX_bit_math_h_l816_c3_7279_iffalse,
layer1_node8_MUX_bit_math_h_l816_c3_7279_return_output);

-- layer1_node9_MUX_bit_math_h_l827_c3_90fc
layer1_node9_MUX_bit_math_h_l827_c3_90fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node9_MUX_bit_math_h_l827_c3_90fc_cond,
layer1_node9_MUX_bit_math_h_l827_c3_90fc_iftrue,
layer1_node9_MUX_bit_math_h_l827_c3_90fc_iffalse,
layer1_node9_MUX_bit_math_h_l827_c3_90fc_return_output);

-- layer1_node10_MUX_bit_math_h_l838_c3_e624
layer1_node10_MUX_bit_math_h_l838_c3_e624 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node10_MUX_bit_math_h_l838_c3_e624_cond,
layer1_node10_MUX_bit_math_h_l838_c3_e624_iftrue,
layer1_node10_MUX_bit_math_h_l838_c3_e624_iffalse,
layer1_node10_MUX_bit_math_h_l838_c3_e624_return_output);

-- layer1_node11_MUX_bit_math_h_l849_c3_0669
layer1_node11_MUX_bit_math_h_l849_c3_0669 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node11_MUX_bit_math_h_l849_c3_0669_cond,
layer1_node11_MUX_bit_math_h_l849_c3_0669_iftrue,
layer1_node11_MUX_bit_math_h_l849_c3_0669_iffalse,
layer1_node11_MUX_bit_math_h_l849_c3_0669_return_output);

-- layer1_node12_MUX_bit_math_h_l860_c3_f017
layer1_node12_MUX_bit_math_h_l860_c3_f017 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node12_MUX_bit_math_h_l860_c3_f017_cond,
layer1_node12_MUX_bit_math_h_l860_c3_f017_iftrue,
layer1_node12_MUX_bit_math_h_l860_c3_f017_iffalse,
layer1_node12_MUX_bit_math_h_l860_c3_f017_return_output);

-- layer1_node13_MUX_bit_math_h_l871_c3_9f0e
layer1_node13_MUX_bit_math_h_l871_c3_9f0e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node13_MUX_bit_math_h_l871_c3_9f0e_cond,
layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iftrue,
layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iffalse,
layer1_node13_MUX_bit_math_h_l871_c3_9f0e_return_output);

-- layer1_node14_MUX_bit_math_h_l882_c3_9be0
layer1_node14_MUX_bit_math_h_l882_c3_9be0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node14_MUX_bit_math_h_l882_c3_9be0_cond,
layer1_node14_MUX_bit_math_h_l882_c3_9be0_iftrue,
layer1_node14_MUX_bit_math_h_l882_c3_9be0_iffalse,
layer1_node14_MUX_bit_math_h_l882_c3_9be0_return_output);

-- layer1_node15_MUX_bit_math_h_l893_c3_db88
layer1_node15_MUX_bit_math_h_l893_c3_db88 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node15_MUX_bit_math_h_l893_c3_db88_cond,
layer1_node15_MUX_bit_math_h_l893_c3_db88_iftrue,
layer1_node15_MUX_bit_math_h_l893_c3_db88_iffalse,
layer1_node15_MUX_bit_math_h_l893_c3_db88_return_output);

-- layer1_node16_MUX_bit_math_h_l904_c3_fdb3
layer1_node16_MUX_bit_math_h_l904_c3_fdb3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node16_MUX_bit_math_h_l904_c3_fdb3_cond,
layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iftrue,
layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iffalse,
layer1_node16_MUX_bit_math_h_l904_c3_fdb3_return_output);

-- layer1_node17_MUX_bit_math_h_l915_c3_bba5
layer1_node17_MUX_bit_math_h_l915_c3_bba5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node17_MUX_bit_math_h_l915_c3_bba5_cond,
layer1_node17_MUX_bit_math_h_l915_c3_bba5_iftrue,
layer1_node17_MUX_bit_math_h_l915_c3_bba5_iffalse,
layer1_node17_MUX_bit_math_h_l915_c3_bba5_return_output);

-- layer1_node18_MUX_bit_math_h_l926_c3_ab1a
layer1_node18_MUX_bit_math_h_l926_c3_ab1a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node18_MUX_bit_math_h_l926_c3_ab1a_cond,
layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iftrue,
layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iffalse,
layer1_node18_MUX_bit_math_h_l926_c3_ab1a_return_output);

-- layer1_node19_MUX_bit_math_h_l937_c3_1a24
layer1_node19_MUX_bit_math_h_l937_c3_1a24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node19_MUX_bit_math_h_l937_c3_1a24_cond,
layer1_node19_MUX_bit_math_h_l937_c3_1a24_iftrue,
layer1_node19_MUX_bit_math_h_l937_c3_1a24_iffalse,
layer1_node19_MUX_bit_math_h_l937_c3_1a24_return_output);

-- layer1_node20_MUX_bit_math_h_l948_c3_2dbc
layer1_node20_MUX_bit_math_h_l948_c3_2dbc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node20_MUX_bit_math_h_l948_c3_2dbc_cond,
layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iftrue,
layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iffalse,
layer1_node20_MUX_bit_math_h_l948_c3_2dbc_return_output);

-- layer1_node21_MUX_bit_math_h_l959_c3_f718
layer1_node21_MUX_bit_math_h_l959_c3_f718 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node21_MUX_bit_math_h_l959_c3_f718_cond,
layer1_node21_MUX_bit_math_h_l959_c3_f718_iftrue,
layer1_node21_MUX_bit_math_h_l959_c3_f718_iffalse,
layer1_node21_MUX_bit_math_h_l959_c3_f718_return_output);

-- layer1_node22_MUX_bit_math_h_l970_c3_3aa5
layer1_node22_MUX_bit_math_h_l970_c3_3aa5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node22_MUX_bit_math_h_l970_c3_3aa5_cond,
layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iftrue,
layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iffalse,
layer1_node22_MUX_bit_math_h_l970_c3_3aa5_return_output);

-- layer1_node23_MUX_bit_math_h_l981_c3_d2b9
layer1_node23_MUX_bit_math_h_l981_c3_d2b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node23_MUX_bit_math_h_l981_c3_d2b9_cond,
layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iftrue,
layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iffalse,
layer1_node23_MUX_bit_math_h_l981_c3_d2b9_return_output);

-- layer1_node24_MUX_bit_math_h_l992_c3_8792
layer1_node24_MUX_bit_math_h_l992_c3_8792 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node24_MUX_bit_math_h_l992_c3_8792_cond,
layer1_node24_MUX_bit_math_h_l992_c3_8792_iftrue,
layer1_node24_MUX_bit_math_h_l992_c3_8792_iffalse,
layer1_node24_MUX_bit_math_h_l992_c3_8792_return_output);

-- layer1_node25_MUX_bit_math_h_l1003_c3_2c90
layer1_node25_MUX_bit_math_h_l1003_c3_2c90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node25_MUX_bit_math_h_l1003_c3_2c90_cond,
layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iftrue,
layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iffalse,
layer1_node25_MUX_bit_math_h_l1003_c3_2c90_return_output);

-- layer1_node26_MUX_bit_math_h_l1014_c3_f8c1
layer1_node26_MUX_bit_math_h_l1014_c3_f8c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_cond,
layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iftrue,
layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iffalse,
layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_return_output);

-- layer1_node27_MUX_bit_math_h_l1025_c3_7ac4
layer1_node27_MUX_bit_math_h_l1025_c3_7ac4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_cond,
layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iftrue,
layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iffalse,
layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_return_output);

-- layer1_node28_MUX_bit_math_h_l1036_c3_deef
layer1_node28_MUX_bit_math_h_l1036_c3_deef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node28_MUX_bit_math_h_l1036_c3_deef_cond,
layer1_node28_MUX_bit_math_h_l1036_c3_deef_iftrue,
layer1_node28_MUX_bit_math_h_l1036_c3_deef_iffalse,
layer1_node28_MUX_bit_math_h_l1036_c3_deef_return_output);

-- layer1_node29_MUX_bit_math_h_l1047_c3_d4d6
layer1_node29_MUX_bit_math_h_l1047_c3_d4d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_cond,
layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iftrue,
layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iffalse,
layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_return_output);

-- layer1_node30_MUX_bit_math_h_l1058_c3_d1f5
layer1_node30_MUX_bit_math_h_l1058_c3_d1f5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_cond,
layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iftrue,
layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iffalse,
layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_return_output);

-- layer1_node31_MUX_bit_math_h_l1069_c3_fc71
layer1_node31_MUX_bit_math_h_l1069_c3_fc71 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node31_MUX_bit_math_h_l1069_c3_fc71_cond,
layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iftrue,
layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iffalse,
layer1_node31_MUX_bit_math_h_l1069_c3_fc71_return_output);

-- layer2_node0_MUX_bit_math_h_l1086_c3_5a52
layer2_node0_MUX_bit_math_h_l1086_c3_5a52 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l1086_c3_5a52_cond,
layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iftrue,
layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iffalse,
layer2_node0_MUX_bit_math_h_l1086_c3_5a52_return_output);

-- layer2_node1_MUX_bit_math_h_l1097_c3_fc1c
layer2_node1_MUX_bit_math_h_l1097_c3_fc1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_cond,
layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iftrue,
layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iffalse,
layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_return_output);

-- layer2_node2_MUX_bit_math_h_l1108_c3_922a
layer2_node2_MUX_bit_math_h_l1108_c3_922a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node2_MUX_bit_math_h_l1108_c3_922a_cond,
layer2_node2_MUX_bit_math_h_l1108_c3_922a_iftrue,
layer2_node2_MUX_bit_math_h_l1108_c3_922a_iffalse,
layer2_node2_MUX_bit_math_h_l1108_c3_922a_return_output);

-- layer2_node3_MUX_bit_math_h_l1119_c3_b25e
layer2_node3_MUX_bit_math_h_l1119_c3_b25e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node3_MUX_bit_math_h_l1119_c3_b25e_cond,
layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iftrue,
layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iffalse,
layer2_node3_MUX_bit_math_h_l1119_c3_b25e_return_output);

-- layer2_node4_MUX_bit_math_h_l1130_c3_5fd5
layer2_node4_MUX_bit_math_h_l1130_c3_5fd5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_cond,
layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iftrue,
layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iffalse,
layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_return_output);

-- layer2_node5_MUX_bit_math_h_l1141_c3_6ecd
layer2_node5_MUX_bit_math_h_l1141_c3_6ecd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_cond,
layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iftrue,
layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iffalse,
layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_return_output);

-- layer2_node6_MUX_bit_math_h_l1152_c3_d917
layer2_node6_MUX_bit_math_h_l1152_c3_d917 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node6_MUX_bit_math_h_l1152_c3_d917_cond,
layer2_node6_MUX_bit_math_h_l1152_c3_d917_iftrue,
layer2_node6_MUX_bit_math_h_l1152_c3_d917_iffalse,
layer2_node6_MUX_bit_math_h_l1152_c3_d917_return_output);

-- layer2_node7_MUX_bit_math_h_l1163_c3_d44d
layer2_node7_MUX_bit_math_h_l1163_c3_d44d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node7_MUX_bit_math_h_l1163_c3_d44d_cond,
layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iftrue,
layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iffalse,
layer2_node7_MUX_bit_math_h_l1163_c3_d44d_return_output);

-- layer2_node8_MUX_bit_math_h_l1174_c3_d504
layer2_node8_MUX_bit_math_h_l1174_c3_d504 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node8_MUX_bit_math_h_l1174_c3_d504_cond,
layer2_node8_MUX_bit_math_h_l1174_c3_d504_iftrue,
layer2_node8_MUX_bit_math_h_l1174_c3_d504_iffalse,
layer2_node8_MUX_bit_math_h_l1174_c3_d504_return_output);

-- layer2_node9_MUX_bit_math_h_l1185_c3_8a90
layer2_node9_MUX_bit_math_h_l1185_c3_8a90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node9_MUX_bit_math_h_l1185_c3_8a90_cond,
layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iftrue,
layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iffalse,
layer2_node9_MUX_bit_math_h_l1185_c3_8a90_return_output);

-- layer2_node10_MUX_bit_math_h_l1196_c3_c6ad
layer2_node10_MUX_bit_math_h_l1196_c3_c6ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_cond,
layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iftrue,
layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iffalse,
layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_return_output);

-- layer2_node11_MUX_bit_math_h_l1207_c3_e593
layer2_node11_MUX_bit_math_h_l1207_c3_e593 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node11_MUX_bit_math_h_l1207_c3_e593_cond,
layer2_node11_MUX_bit_math_h_l1207_c3_e593_iftrue,
layer2_node11_MUX_bit_math_h_l1207_c3_e593_iffalse,
layer2_node11_MUX_bit_math_h_l1207_c3_e593_return_output);

-- layer2_node12_MUX_bit_math_h_l1218_c3_ed0c
layer2_node12_MUX_bit_math_h_l1218_c3_ed0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_cond,
layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iftrue,
layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iffalse,
layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_return_output);

-- layer2_node13_MUX_bit_math_h_l1229_c3_d88d
layer2_node13_MUX_bit_math_h_l1229_c3_d88d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node13_MUX_bit_math_h_l1229_c3_d88d_cond,
layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iftrue,
layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iffalse,
layer2_node13_MUX_bit_math_h_l1229_c3_d88d_return_output);

-- layer2_node14_MUX_bit_math_h_l1240_c3_d3d6
layer2_node14_MUX_bit_math_h_l1240_c3_d3d6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_cond,
layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iftrue,
layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iffalse,
layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_return_output);

-- layer2_node15_MUX_bit_math_h_l1251_c3_03ac
layer2_node15_MUX_bit_math_h_l1251_c3_03ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node15_MUX_bit_math_h_l1251_c3_03ac_cond,
layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iftrue,
layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iffalse,
layer2_node15_MUX_bit_math_h_l1251_c3_03ac_return_output);

-- layer3_node0_MUX_bit_math_h_l1268_c3_6917
layer3_node0_MUX_bit_math_h_l1268_c3_6917 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l1268_c3_6917_cond,
layer3_node0_MUX_bit_math_h_l1268_c3_6917_iftrue,
layer3_node0_MUX_bit_math_h_l1268_c3_6917_iffalse,
layer3_node0_MUX_bit_math_h_l1268_c3_6917_return_output);

-- layer3_node1_MUX_bit_math_h_l1279_c3_e270
layer3_node1_MUX_bit_math_h_l1279_c3_e270 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node1_MUX_bit_math_h_l1279_c3_e270_cond,
layer3_node1_MUX_bit_math_h_l1279_c3_e270_iftrue,
layer3_node1_MUX_bit_math_h_l1279_c3_e270_iffalse,
layer3_node1_MUX_bit_math_h_l1279_c3_e270_return_output);

-- layer3_node2_MUX_bit_math_h_l1290_c3_769c
layer3_node2_MUX_bit_math_h_l1290_c3_769c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node2_MUX_bit_math_h_l1290_c3_769c_cond,
layer3_node2_MUX_bit_math_h_l1290_c3_769c_iftrue,
layer3_node2_MUX_bit_math_h_l1290_c3_769c_iffalse,
layer3_node2_MUX_bit_math_h_l1290_c3_769c_return_output);

-- layer3_node3_MUX_bit_math_h_l1301_c3_fb21
layer3_node3_MUX_bit_math_h_l1301_c3_fb21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node3_MUX_bit_math_h_l1301_c3_fb21_cond,
layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iftrue,
layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iffalse,
layer3_node3_MUX_bit_math_h_l1301_c3_fb21_return_output);

-- layer3_node4_MUX_bit_math_h_l1312_c3_f274
layer3_node4_MUX_bit_math_h_l1312_c3_f274 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node4_MUX_bit_math_h_l1312_c3_f274_cond,
layer3_node4_MUX_bit_math_h_l1312_c3_f274_iftrue,
layer3_node4_MUX_bit_math_h_l1312_c3_f274_iffalse,
layer3_node4_MUX_bit_math_h_l1312_c3_f274_return_output);

-- layer3_node5_MUX_bit_math_h_l1323_c3_6b46
layer3_node5_MUX_bit_math_h_l1323_c3_6b46 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node5_MUX_bit_math_h_l1323_c3_6b46_cond,
layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iftrue,
layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iffalse,
layer3_node5_MUX_bit_math_h_l1323_c3_6b46_return_output);

-- layer3_node6_MUX_bit_math_h_l1334_c3_41a0
layer3_node6_MUX_bit_math_h_l1334_c3_41a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node6_MUX_bit_math_h_l1334_c3_41a0_cond,
layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iftrue,
layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iffalse,
layer3_node6_MUX_bit_math_h_l1334_c3_41a0_return_output);

-- layer3_node7_MUX_bit_math_h_l1345_c3_969c
layer3_node7_MUX_bit_math_h_l1345_c3_969c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node7_MUX_bit_math_h_l1345_c3_969c_cond,
layer3_node7_MUX_bit_math_h_l1345_c3_969c_iftrue,
layer3_node7_MUX_bit_math_h_l1345_c3_969c_iffalse,
layer3_node7_MUX_bit_math_h_l1345_c3_969c_return_output);

-- layer4_node0_MUX_bit_math_h_l1362_c3_b41d
layer4_node0_MUX_bit_math_h_l1362_c3_b41d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node0_MUX_bit_math_h_l1362_c3_b41d_cond,
layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iftrue,
layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iffalse,
layer4_node0_MUX_bit_math_h_l1362_c3_b41d_return_output);

-- layer4_node1_MUX_bit_math_h_l1373_c3_f2a6
layer4_node1_MUX_bit_math_h_l1373_c3_f2a6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_cond,
layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iftrue,
layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iffalse,
layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_return_output);

-- layer4_node2_MUX_bit_math_h_l1384_c3_3339
layer4_node2_MUX_bit_math_h_l1384_c3_3339 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node2_MUX_bit_math_h_l1384_c3_3339_cond,
layer4_node2_MUX_bit_math_h_l1384_c3_3339_iftrue,
layer4_node2_MUX_bit_math_h_l1384_c3_3339_iffalse,
layer4_node2_MUX_bit_math_h_l1384_c3_3339_return_output);

-- layer4_node3_MUX_bit_math_h_l1395_c3_b75d
layer4_node3_MUX_bit_math_h_l1395_c3_b75d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node3_MUX_bit_math_h_l1395_c3_b75d_cond,
layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iftrue,
layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iffalse,
layer4_node3_MUX_bit_math_h_l1395_c3_b75d_return_output);

-- layer5_node0_MUX_bit_math_h_l1412_c3_5f1f
layer5_node0_MUX_bit_math_h_l1412_c3_5f1f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_cond,
layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iftrue,
layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iffalse,
layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_return_output);

-- layer5_node1_MUX_bit_math_h_l1423_c3_1d22
layer5_node1_MUX_bit_math_h_l1423_c3_1d22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node1_MUX_bit_math_h_l1423_c3_1d22_cond,
layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iftrue,
layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iffalse,
layer5_node1_MUX_bit_math_h_l1423_c3_1d22_return_output);

-- layer6_node0_MUX_bit_math_h_l1440_c3_247e
layer6_node0_MUX_bit_math_h_l1440_c3_247e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer6_node0_MUX_bit_math_h_l1440_c3_247e_cond,
layer6_node0_MUX_bit_math_h_l1440_c3_247e_iftrue,
layer6_node0_MUX_bit_math_h_l1440_c3_247e_iffalse,
layer6_node0_MUX_bit_math_h_l1440_c3_247e_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 in16,
 in17,
 in18,
 in19,
 in20,
 in21,
 in22,
 in23,
 in24,
 in25,
 in26,
 in27,
 in28,
 in29,
 in30,
 in31,
 in32,
 in33,
 in34,
 in35,
 in36,
 in37,
 in38,
 in39,
 in40,
 in41,
 in42,
 in43,
 in44,
 in45,
 in46,
 in47,
 in48,
 in49,
 in50,
 in51,
 in52,
 in53,
 in54,
 in55,
 in56,
 in57,
 in58,
 in59,
 in60,
 in61,
 in62,
 in63,
 in64,
 in65,
 in66,
 in67,
 in68,
 in69,
 in70,
 in71,
 in72,
 in73,
 in74,
 in75,
 in76,
 in77,
 in78,
 in79,
 in80,
 in81,
 in82,
 in83,
 in84,
 in85,
 in86,
 in87,
 in88,
 in89,
 in90,
 in91,
 in92,
 in93,
 in94,
 in95,
 in96,
 in97,
 in98,
 in99,
 in100,
 in101,
 in102,
 in103,
 in104,
 in105,
 in106,
 in107,
 in108,
 in109,
 in110,
 in111,
 in112,
 in113,
 in114,
 in115,
 in116,
 in117,
 in118,
 in119,
 in120,
 in121,
 in122,
 in123,
 in124,
 in125,
 in126,
 in127,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_8bd4_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_b2fc_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_3d12_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_13b9_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_be4c_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_936b_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_6f9a_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_f259_return_output,
 layer0_node8_MUX_bit_math_h_l106_c3_2e0c_return_output,
 layer0_node9_MUX_bit_math_h_l117_c3_1a47_return_output,
 layer0_node10_MUX_bit_math_h_l128_c3_0e40_return_output,
 layer0_node11_MUX_bit_math_h_l139_c3_381c_return_output,
 layer0_node12_MUX_bit_math_h_l150_c3_1560_return_output,
 layer0_node13_MUX_bit_math_h_l161_c3_3a1c_return_output,
 layer0_node14_MUX_bit_math_h_l172_c3_7ef7_return_output,
 layer0_node15_MUX_bit_math_h_l183_c3_392b_return_output,
 layer0_node16_MUX_bit_math_h_l194_c3_cada_return_output,
 layer0_node17_MUX_bit_math_h_l205_c3_39fd_return_output,
 layer0_node18_MUX_bit_math_h_l216_c3_23c8_return_output,
 layer0_node19_MUX_bit_math_h_l227_c3_ea58_return_output,
 layer0_node20_MUX_bit_math_h_l238_c3_eb78_return_output,
 layer0_node21_MUX_bit_math_h_l249_c3_228d_return_output,
 layer0_node22_MUX_bit_math_h_l260_c3_1c3c_return_output,
 layer0_node23_MUX_bit_math_h_l271_c3_6340_return_output,
 layer0_node24_MUX_bit_math_h_l282_c3_670b_return_output,
 layer0_node25_MUX_bit_math_h_l293_c3_83e8_return_output,
 layer0_node26_MUX_bit_math_h_l304_c3_53e2_return_output,
 layer0_node27_MUX_bit_math_h_l315_c3_ac24_return_output,
 layer0_node28_MUX_bit_math_h_l326_c3_97ed_return_output,
 layer0_node29_MUX_bit_math_h_l337_c3_7a23_return_output,
 layer0_node30_MUX_bit_math_h_l348_c3_7ed3_return_output,
 layer0_node31_MUX_bit_math_h_l359_c3_208c_return_output,
 layer0_node32_MUX_bit_math_h_l370_c3_bcd8_return_output,
 layer0_node33_MUX_bit_math_h_l381_c3_0aac_return_output,
 layer0_node34_MUX_bit_math_h_l392_c3_6801_return_output,
 layer0_node35_MUX_bit_math_h_l403_c3_749b_return_output,
 layer0_node36_MUX_bit_math_h_l414_c3_0db7_return_output,
 layer0_node37_MUX_bit_math_h_l425_c3_7f65_return_output,
 layer0_node38_MUX_bit_math_h_l436_c3_d774_return_output,
 layer0_node39_MUX_bit_math_h_l447_c3_b0c4_return_output,
 layer0_node40_MUX_bit_math_h_l458_c3_773e_return_output,
 layer0_node41_MUX_bit_math_h_l469_c3_62cc_return_output,
 layer0_node42_MUX_bit_math_h_l480_c3_d626_return_output,
 layer0_node43_MUX_bit_math_h_l491_c3_001b_return_output,
 layer0_node44_MUX_bit_math_h_l502_c3_1816_return_output,
 layer0_node45_MUX_bit_math_h_l513_c3_cc83_return_output,
 layer0_node46_MUX_bit_math_h_l524_c3_aa0a_return_output,
 layer0_node47_MUX_bit_math_h_l535_c3_167a_return_output,
 layer0_node48_MUX_bit_math_h_l546_c3_41a2_return_output,
 layer0_node49_MUX_bit_math_h_l557_c3_3c6d_return_output,
 layer0_node50_MUX_bit_math_h_l568_c3_e0e2_return_output,
 layer0_node51_MUX_bit_math_h_l579_c3_1b2f_return_output,
 layer0_node52_MUX_bit_math_h_l590_c3_dee1_return_output,
 layer0_node53_MUX_bit_math_h_l601_c3_76ac_return_output,
 layer0_node54_MUX_bit_math_h_l612_c3_e1c8_return_output,
 layer0_node55_MUX_bit_math_h_l623_c3_ec7e_return_output,
 layer0_node56_MUX_bit_math_h_l634_c3_5b10_return_output,
 layer0_node57_MUX_bit_math_h_l645_c3_d7f5_return_output,
 layer0_node58_MUX_bit_math_h_l656_c3_e8c0_return_output,
 layer0_node59_MUX_bit_math_h_l667_c3_1ea2_return_output,
 layer0_node60_MUX_bit_math_h_l678_c3_fe9f_return_output,
 layer0_node61_MUX_bit_math_h_l689_c3_9f98_return_output,
 layer0_node62_MUX_bit_math_h_l700_c3_0d13_return_output,
 layer0_node63_MUX_bit_math_h_l711_c3_2778_return_output,
 layer1_node0_MUX_bit_math_h_l728_c3_67cd_return_output,
 layer1_node1_MUX_bit_math_h_l739_c3_5e54_return_output,
 layer1_node2_MUX_bit_math_h_l750_c3_386d_return_output,
 layer1_node3_MUX_bit_math_h_l761_c3_c96d_return_output,
 layer1_node4_MUX_bit_math_h_l772_c3_535b_return_output,
 layer1_node5_MUX_bit_math_h_l783_c3_7132_return_output,
 layer1_node6_MUX_bit_math_h_l794_c3_59a7_return_output,
 layer1_node7_MUX_bit_math_h_l805_c3_a7b7_return_output,
 layer1_node8_MUX_bit_math_h_l816_c3_7279_return_output,
 layer1_node9_MUX_bit_math_h_l827_c3_90fc_return_output,
 layer1_node10_MUX_bit_math_h_l838_c3_e624_return_output,
 layer1_node11_MUX_bit_math_h_l849_c3_0669_return_output,
 layer1_node12_MUX_bit_math_h_l860_c3_f017_return_output,
 layer1_node13_MUX_bit_math_h_l871_c3_9f0e_return_output,
 layer1_node14_MUX_bit_math_h_l882_c3_9be0_return_output,
 layer1_node15_MUX_bit_math_h_l893_c3_db88_return_output,
 layer1_node16_MUX_bit_math_h_l904_c3_fdb3_return_output,
 layer1_node17_MUX_bit_math_h_l915_c3_bba5_return_output,
 layer1_node18_MUX_bit_math_h_l926_c3_ab1a_return_output,
 layer1_node19_MUX_bit_math_h_l937_c3_1a24_return_output,
 layer1_node20_MUX_bit_math_h_l948_c3_2dbc_return_output,
 layer1_node21_MUX_bit_math_h_l959_c3_f718_return_output,
 layer1_node22_MUX_bit_math_h_l970_c3_3aa5_return_output,
 layer1_node23_MUX_bit_math_h_l981_c3_d2b9_return_output,
 layer1_node24_MUX_bit_math_h_l992_c3_8792_return_output,
 layer1_node25_MUX_bit_math_h_l1003_c3_2c90_return_output,
 layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_return_output,
 layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_return_output,
 layer1_node28_MUX_bit_math_h_l1036_c3_deef_return_output,
 layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_return_output,
 layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_return_output,
 layer1_node31_MUX_bit_math_h_l1069_c3_fc71_return_output,
 layer2_node0_MUX_bit_math_h_l1086_c3_5a52_return_output,
 layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_return_output,
 layer2_node2_MUX_bit_math_h_l1108_c3_922a_return_output,
 layer2_node3_MUX_bit_math_h_l1119_c3_b25e_return_output,
 layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_return_output,
 layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_return_output,
 layer2_node6_MUX_bit_math_h_l1152_c3_d917_return_output,
 layer2_node7_MUX_bit_math_h_l1163_c3_d44d_return_output,
 layer2_node8_MUX_bit_math_h_l1174_c3_d504_return_output,
 layer2_node9_MUX_bit_math_h_l1185_c3_8a90_return_output,
 layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_return_output,
 layer2_node11_MUX_bit_math_h_l1207_c3_e593_return_output,
 layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_return_output,
 layer2_node13_MUX_bit_math_h_l1229_c3_d88d_return_output,
 layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_return_output,
 layer2_node15_MUX_bit_math_h_l1251_c3_03ac_return_output,
 layer3_node0_MUX_bit_math_h_l1268_c3_6917_return_output,
 layer3_node1_MUX_bit_math_h_l1279_c3_e270_return_output,
 layer3_node2_MUX_bit_math_h_l1290_c3_769c_return_output,
 layer3_node3_MUX_bit_math_h_l1301_c3_fb21_return_output,
 layer3_node4_MUX_bit_math_h_l1312_c3_f274_return_output,
 layer3_node5_MUX_bit_math_h_l1323_c3_6b46_return_output,
 layer3_node6_MUX_bit_math_h_l1334_c3_41a0_return_output,
 layer3_node7_MUX_bit_math_h_l1345_c3_969c_return_output,
 layer4_node0_MUX_bit_math_h_l1362_c3_b41d_return_output,
 layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_return_output,
 layer4_node2_MUX_bit_math_h_l1384_c3_3339_return_output,
 layer4_node3_MUX_bit_math_h_l1395_c3_b75d_return_output,
 layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_return_output,
 layer5_node1_MUX_bit_math_h_l1423_c3_1d22_return_output,
 layer6_node0_MUX_bit_math_h_l1440_c3_247e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(7 downto 0);
 variable VAR_sel : unsigned(6 downto 0);
 variable VAR_in0 : unsigned(7 downto 0);
 variable VAR_in1 : unsigned(7 downto 0);
 variable VAR_in2 : unsigned(7 downto 0);
 variable VAR_in3 : unsigned(7 downto 0);
 variable VAR_in4 : unsigned(7 downto 0);
 variable VAR_in5 : unsigned(7 downto 0);
 variable VAR_in6 : unsigned(7 downto 0);
 variable VAR_in7 : unsigned(7 downto 0);
 variable VAR_in8 : unsigned(7 downto 0);
 variable VAR_in9 : unsigned(7 downto 0);
 variable VAR_in10 : unsigned(7 downto 0);
 variable VAR_in11 : unsigned(7 downto 0);
 variable VAR_in12 : unsigned(7 downto 0);
 variable VAR_in13 : unsigned(7 downto 0);
 variable VAR_in14 : unsigned(7 downto 0);
 variable VAR_in15 : unsigned(7 downto 0);
 variable VAR_in16 : unsigned(7 downto 0);
 variable VAR_in17 : unsigned(7 downto 0);
 variable VAR_in18 : unsigned(7 downto 0);
 variable VAR_in19 : unsigned(7 downto 0);
 variable VAR_in20 : unsigned(7 downto 0);
 variable VAR_in21 : unsigned(7 downto 0);
 variable VAR_in22 : unsigned(7 downto 0);
 variable VAR_in23 : unsigned(7 downto 0);
 variable VAR_in24 : unsigned(7 downto 0);
 variable VAR_in25 : unsigned(7 downto 0);
 variable VAR_in26 : unsigned(7 downto 0);
 variable VAR_in27 : unsigned(7 downto 0);
 variable VAR_in28 : unsigned(7 downto 0);
 variable VAR_in29 : unsigned(7 downto 0);
 variable VAR_in30 : unsigned(7 downto 0);
 variable VAR_in31 : unsigned(7 downto 0);
 variable VAR_in32 : unsigned(7 downto 0);
 variable VAR_in33 : unsigned(7 downto 0);
 variable VAR_in34 : unsigned(7 downto 0);
 variable VAR_in35 : unsigned(7 downto 0);
 variable VAR_in36 : unsigned(7 downto 0);
 variable VAR_in37 : unsigned(7 downto 0);
 variable VAR_in38 : unsigned(7 downto 0);
 variable VAR_in39 : unsigned(7 downto 0);
 variable VAR_in40 : unsigned(7 downto 0);
 variable VAR_in41 : unsigned(7 downto 0);
 variable VAR_in42 : unsigned(7 downto 0);
 variable VAR_in43 : unsigned(7 downto 0);
 variable VAR_in44 : unsigned(7 downto 0);
 variable VAR_in45 : unsigned(7 downto 0);
 variable VAR_in46 : unsigned(7 downto 0);
 variable VAR_in47 : unsigned(7 downto 0);
 variable VAR_in48 : unsigned(7 downto 0);
 variable VAR_in49 : unsigned(7 downto 0);
 variable VAR_in50 : unsigned(7 downto 0);
 variable VAR_in51 : unsigned(7 downto 0);
 variable VAR_in52 : unsigned(7 downto 0);
 variable VAR_in53 : unsigned(7 downto 0);
 variable VAR_in54 : unsigned(7 downto 0);
 variable VAR_in55 : unsigned(7 downto 0);
 variable VAR_in56 : unsigned(7 downto 0);
 variable VAR_in57 : unsigned(7 downto 0);
 variable VAR_in58 : unsigned(7 downto 0);
 variable VAR_in59 : unsigned(7 downto 0);
 variable VAR_in60 : unsigned(7 downto 0);
 variable VAR_in61 : unsigned(7 downto 0);
 variable VAR_in62 : unsigned(7 downto 0);
 variable VAR_in63 : unsigned(7 downto 0);
 variable VAR_in64 : unsigned(7 downto 0);
 variable VAR_in65 : unsigned(7 downto 0);
 variable VAR_in66 : unsigned(7 downto 0);
 variable VAR_in67 : unsigned(7 downto 0);
 variable VAR_in68 : unsigned(7 downto 0);
 variable VAR_in69 : unsigned(7 downto 0);
 variable VAR_in70 : unsigned(7 downto 0);
 variable VAR_in71 : unsigned(7 downto 0);
 variable VAR_in72 : unsigned(7 downto 0);
 variable VAR_in73 : unsigned(7 downto 0);
 variable VAR_in74 : unsigned(7 downto 0);
 variable VAR_in75 : unsigned(7 downto 0);
 variable VAR_in76 : unsigned(7 downto 0);
 variable VAR_in77 : unsigned(7 downto 0);
 variable VAR_in78 : unsigned(7 downto 0);
 variable VAR_in79 : unsigned(7 downto 0);
 variable VAR_in80 : unsigned(7 downto 0);
 variable VAR_in81 : unsigned(7 downto 0);
 variable VAR_in82 : unsigned(7 downto 0);
 variable VAR_in83 : unsigned(7 downto 0);
 variable VAR_in84 : unsigned(7 downto 0);
 variable VAR_in85 : unsigned(7 downto 0);
 variable VAR_in86 : unsigned(7 downto 0);
 variable VAR_in87 : unsigned(7 downto 0);
 variable VAR_in88 : unsigned(7 downto 0);
 variable VAR_in89 : unsigned(7 downto 0);
 variable VAR_in90 : unsigned(7 downto 0);
 variable VAR_in91 : unsigned(7 downto 0);
 variable VAR_in92 : unsigned(7 downto 0);
 variable VAR_in93 : unsigned(7 downto 0);
 variable VAR_in94 : unsigned(7 downto 0);
 variable VAR_in95 : unsigned(7 downto 0);
 variable VAR_in96 : unsigned(7 downto 0);
 variable VAR_in97 : unsigned(7 downto 0);
 variable VAR_in98 : unsigned(7 downto 0);
 variable VAR_in99 : unsigned(7 downto 0);
 variable VAR_in100 : unsigned(7 downto 0);
 variable VAR_in101 : unsigned(7 downto 0);
 variable VAR_in102 : unsigned(7 downto 0);
 variable VAR_in103 : unsigned(7 downto 0);
 variable VAR_in104 : unsigned(7 downto 0);
 variable VAR_in105 : unsigned(7 downto 0);
 variable VAR_in106 : unsigned(7 downto 0);
 variable VAR_in107 : unsigned(7 downto 0);
 variable VAR_in108 : unsigned(7 downto 0);
 variable VAR_in109 : unsigned(7 downto 0);
 variable VAR_in110 : unsigned(7 downto 0);
 variable VAR_in111 : unsigned(7 downto 0);
 variable VAR_in112 : unsigned(7 downto 0);
 variable VAR_in113 : unsigned(7 downto 0);
 variable VAR_in114 : unsigned(7 downto 0);
 variable VAR_in115 : unsigned(7 downto 0);
 variable VAR_in116 : unsigned(7 downto 0);
 variable VAR_in117 : unsigned(7 downto 0);
 variable VAR_in118 : unsigned(7 downto 0);
 variable VAR_in119 : unsigned(7 downto 0);
 variable VAR_in120 : unsigned(7 downto 0);
 variable VAR_in121 : unsigned(7 downto 0);
 variable VAR_in122 : unsigned(7 downto 0);
 variable VAR_in123 : unsigned(7 downto 0);
 variable VAR_in124 : unsigned(7 downto 0);
 variable VAR_in125 : unsigned(7 downto 0);
 variable VAR_in126 : unsigned(7 downto 0);
 variable VAR_in127 : unsigned(7 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_cond : unsigned(0 downto 0);
 variable VAR_layer0_node8 : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node9 : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_cond : unsigned(0 downto 0);
 variable VAR_layer0_node10 : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_cond : unsigned(0 downto 0);
 variable VAR_layer0_node11 : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node12 : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_cond : unsigned(0 downto 0);
 variable VAR_layer0_node13 : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node14 : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node15 : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node16 : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_cond : unsigned(0 downto 0);
 variable VAR_layer0_node17 : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_cond : unsigned(0 downto 0);
 variable VAR_layer0_node18 : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node19 : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_cond : unsigned(0 downto 0);
 variable VAR_layer0_node20 : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_cond : unsigned(0 downto 0);
 variable VAR_layer0_node21 : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node22 : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node23 : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_cond : unsigned(0 downto 0);
 variable VAR_layer0_node24 : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node25 : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node26 : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node27 : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_cond : unsigned(0 downto 0);
 variable VAR_layer0_node28 : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_cond : unsigned(0 downto 0);
 variable VAR_layer0_node29 : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_cond : unsigned(0 downto 0);
 variable VAR_layer0_node30 : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node31 : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node32 : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node33 : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_cond : unsigned(0 downto 0);
 variable VAR_layer0_node34 : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_cond : unsigned(0 downto 0);
 variable VAR_layer0_node35 : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node36 : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node37 : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_cond : unsigned(0 downto 0);
 variable VAR_layer0_node38 : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_cond : unsigned(0 downto 0);
 variable VAR_layer0_node39 : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_cond : unsigned(0 downto 0);
 variable VAR_layer0_node40 : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node41 : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_cond : unsigned(0 downto 0);
 variable VAR_layer0_node42 : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_cond : unsigned(0 downto 0);
 variable VAR_layer0_node43 : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node44 : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_cond : unsigned(0 downto 0);
 variable VAR_layer0_node45 : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_cond : unsigned(0 downto 0);
 variable VAR_layer0_node46 : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node47 : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node48 : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node49 : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node50 : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node51 : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_cond : unsigned(0 downto 0);
 variable VAR_layer0_node52 : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node53 : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_cond : unsigned(0 downto 0);
 variable VAR_layer0_node54 : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node55 : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node56 : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_cond : unsigned(0 downto 0);
 variable VAR_layer0_node57 : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_cond : unsigned(0 downto 0);
 variable VAR_layer0_node58 : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_cond : unsigned(0 downto 0);
 variable VAR_layer0_node59 : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_cond : unsigned(0 downto 0);
 variable VAR_layer0_node60 : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_cond : unsigned(0 downto 0);
 variable VAR_layer0_node61 : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_cond : unsigned(0 downto 0);
 variable VAR_layer0_node62 : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_cond : unsigned(0 downto 0);
 variable VAR_layer0_node63 : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_cond : unsigned(0 downto 0);
 variable VAR_layer1_node4 : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_cond : unsigned(0 downto 0);
 variable VAR_layer1_node5 : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_cond : unsigned(0 downto 0);
 variable VAR_layer1_node6 : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_cond : unsigned(0 downto 0);
 variable VAR_layer1_node7 : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_cond : unsigned(0 downto 0);
 variable VAR_layer1_node8 : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_cond : unsigned(0 downto 0);
 variable VAR_layer1_node9 : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_cond : unsigned(0 downto 0);
 variable VAR_layer1_node10 : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_cond : unsigned(0 downto 0);
 variable VAR_layer1_node11 : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_cond : unsigned(0 downto 0);
 variable VAR_layer1_node12 : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_cond : unsigned(0 downto 0);
 variable VAR_layer1_node13 : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_cond : unsigned(0 downto 0);
 variable VAR_layer1_node14 : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_cond : unsigned(0 downto 0);
 variable VAR_layer1_node15 : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_cond : unsigned(0 downto 0);
 variable VAR_layer1_node16 : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_cond : unsigned(0 downto 0);
 variable VAR_layer1_node17 : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_cond : unsigned(0 downto 0);
 variable VAR_layer1_node18 : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_cond : unsigned(0 downto 0);
 variable VAR_layer1_node19 : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_cond : unsigned(0 downto 0);
 variable VAR_layer1_node20 : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_cond : unsigned(0 downto 0);
 variable VAR_layer1_node21 : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_cond : unsigned(0 downto 0);
 variable VAR_layer1_node22 : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_cond : unsigned(0 downto 0);
 variable VAR_layer1_node23 : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_cond : unsigned(0 downto 0);
 variable VAR_layer1_node24 : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_cond : unsigned(0 downto 0);
 variable VAR_layer1_node25 : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_cond : unsigned(0 downto 0);
 variable VAR_layer1_node26 : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_cond : unsigned(0 downto 0);
 variable VAR_layer1_node27 : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_cond : unsigned(0 downto 0);
 variable VAR_layer1_node28 : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_cond : unsigned(0 downto 0);
 variable VAR_layer1_node29 : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_cond : unsigned(0 downto 0);
 variable VAR_layer1_node30 : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_cond : unsigned(0 downto 0);
 variable VAR_layer1_node31 : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_cond : unsigned(0 downto 0);
 variable VAR_layer2_node2 : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_cond : unsigned(0 downto 0);
 variable VAR_layer2_node3 : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_cond : unsigned(0 downto 0);
 variable VAR_layer2_node4 : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_cond : unsigned(0 downto 0);
 variable VAR_layer2_node5 : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_cond : unsigned(0 downto 0);
 variable VAR_layer2_node6 : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_cond : unsigned(0 downto 0);
 variable VAR_layer2_node7 : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_cond : unsigned(0 downto 0);
 variable VAR_layer2_node8 : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_cond : unsigned(0 downto 0);
 variable VAR_layer2_node9 : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_cond : unsigned(0 downto 0);
 variable VAR_layer2_node10 : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_cond : unsigned(0 downto 0);
 variable VAR_layer2_node11 : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_cond : unsigned(0 downto 0);
 variable VAR_layer2_node12 : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_cond : unsigned(0 downto 0);
 variable VAR_layer2_node13 : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_cond : unsigned(0 downto 0);
 variable VAR_layer2_node14 : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_cond : unsigned(0 downto 0);
 variable VAR_layer2_node15 : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_cond : unsigned(0 downto 0);
 variable VAR_layer3_node1 : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_cond : unsigned(0 downto 0);
 variable VAR_layer3_node2 : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_cond : unsigned(0 downto 0);
 variable VAR_layer3_node3 : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_cond : unsigned(0 downto 0);
 variable VAR_layer3_node4 : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_cond : unsigned(0 downto 0);
 variable VAR_layer3_node5 : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_cond : unsigned(0 downto 0);
 variable VAR_layer3_node6 : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_cond : unsigned(0 downto 0);
 variable VAR_layer3_node7 : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_cond : unsigned(0 downto 0);
 variable VAR_sel4 : unsigned(0 downto 0);
 variable VAR_uint7_4_4_bit_math_h_l1358_c10_c24c_return_output : unsigned(0 downto 0);
 variable VAR_layer4_node0 : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_cond : unsigned(0 downto 0);
 variable VAR_layer4_node1 : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_cond : unsigned(0 downto 0);
 variable VAR_layer4_node2 : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_cond : unsigned(0 downto 0);
 variable VAR_layer4_node3 : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_cond : unsigned(0 downto 0);
 variable VAR_sel5 : unsigned(0 downto 0);
 variable VAR_uint7_5_5_bit_math_h_l1408_c10_901f_return_output : unsigned(0 downto 0);
 variable VAR_layer5_node0 : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_cond : unsigned(0 downto 0);
 variable VAR_layer5_node1 : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_cond : unsigned(0 downto 0);
 variable VAR_sel6 : unsigned(0 downto 0);
 variable VAR_uint7_6_6_bit_math_h_l1436_c10_87f9_return_output : unsigned(0 downto 0);
 variable VAR_layer6_node0 : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_iftrue : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_iffalse : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_return_output : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;
     VAR_in16 := in16;
     VAR_in17 := in17;
     VAR_in18 := in18;
     VAR_in19 := in19;
     VAR_in20 := in20;
     VAR_in21 := in21;
     VAR_in22 := in22;
     VAR_in23 := in23;
     VAR_in24 := in24;
     VAR_in25 := in25;
     VAR_in26 := in26;
     VAR_in27 := in27;
     VAR_in28 := in28;
     VAR_in29 := in29;
     VAR_in30 := in30;
     VAR_in31 := in31;
     VAR_in32 := in32;
     VAR_in33 := in33;
     VAR_in34 := in34;
     VAR_in35 := in35;
     VAR_in36 := in36;
     VAR_in37 := in37;
     VAR_in38 := in38;
     VAR_in39 := in39;
     VAR_in40 := in40;
     VAR_in41 := in41;
     VAR_in42 := in42;
     VAR_in43 := in43;
     VAR_in44 := in44;
     VAR_in45 := in45;
     VAR_in46 := in46;
     VAR_in47 := in47;
     VAR_in48 := in48;
     VAR_in49 := in49;
     VAR_in50 := in50;
     VAR_in51 := in51;
     VAR_in52 := in52;
     VAR_in53 := in53;
     VAR_in54 := in54;
     VAR_in55 := in55;
     VAR_in56 := in56;
     VAR_in57 := in57;
     VAR_in58 := in58;
     VAR_in59 := in59;
     VAR_in60 := in60;
     VAR_in61 := in61;
     VAR_in62 := in62;
     VAR_in63 := in63;
     VAR_in64 := in64;
     VAR_in65 := in65;
     VAR_in66 := in66;
     VAR_in67 := in67;
     VAR_in68 := in68;
     VAR_in69 := in69;
     VAR_in70 := in70;
     VAR_in71 := in71;
     VAR_in72 := in72;
     VAR_in73 := in73;
     VAR_in74 := in74;
     VAR_in75 := in75;
     VAR_in76 := in76;
     VAR_in77 := in77;
     VAR_in78 := in78;
     VAR_in79 := in79;
     VAR_in80 := in80;
     VAR_in81 := in81;
     VAR_in82 := in82;
     VAR_in83 := in83;
     VAR_in84 := in84;
     VAR_in85 := in85;
     VAR_in86 := in86;
     VAR_in87 := in87;
     VAR_in88 := in88;
     VAR_in89 := in89;
     VAR_in90 := in90;
     VAR_in91 := in91;
     VAR_in92 := in92;
     VAR_in93 := in93;
     VAR_in94 := in94;
     VAR_in95 := in95;
     VAR_in96 := in96;
     VAR_in97 := in97;
     VAR_in98 := in98;
     VAR_in99 := in99;
     VAR_in100 := in100;
     VAR_in101 := in101;
     VAR_in102 := in102;
     VAR_in103 := in103;
     VAR_in104 := in104;
     VAR_in105 := in105;
     VAR_in106 := in106;
     VAR_in107 := in107;
     VAR_in108 := in108;
     VAR_in109 := in109;
     VAR_in110 := in110;
     VAR_in111 := in111;
     VAR_in112 := in112;
     VAR_in113 := in113;
     VAR_in114 := in114;
     VAR_in115 := in115;
     VAR_in116 := in116;
     VAR_in117 := in117;
     VAR_in118 := in118;
     VAR_in119 := in119;
     VAR_in120 := in120;
     VAR_in121 := in121;
     VAR_in122 := in122;
     VAR_in123 := in123;
     VAR_in124 := in124;
     VAR_in125 := in125;
     VAR_in126 := in126;
     VAR_in127 := in127;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_iffalse := VAR_in10;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iffalse := VAR_in100;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iftrue := VAR_in101;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iffalse := VAR_in102;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iftrue := VAR_in103;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_iffalse := VAR_in104;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_iftrue := VAR_in105;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_iffalse := VAR_in106;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_iftrue := VAR_in107;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iffalse := VAR_in108;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iftrue := VAR_in109;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_iftrue := VAR_in11;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iffalse := VAR_in110;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iftrue := VAR_in111;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_iffalse := VAR_in112;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_iftrue := VAR_in113;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iffalse := VAR_in114;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iftrue := VAR_in115;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iffalse := VAR_in116;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iftrue := VAR_in117;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iffalse := VAR_in118;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iftrue := VAR_in119;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iffalse := VAR_in12;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iffalse := VAR_in120;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iftrue := VAR_in121;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_iffalse := VAR_in122;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_iftrue := VAR_in123;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_iffalse := VAR_in124;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_iftrue := VAR_in125;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_iffalse := VAR_in126;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_iftrue := VAR_in127;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_iftrue := VAR_in15;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iffalse := VAR_in16;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iftrue := VAR_in17;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_iffalse := VAR_in18;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_iftrue := VAR_in19;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iffalse := VAR_in2;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_iffalse := VAR_in20;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_iftrue := VAR_in21;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_iffalse := VAR_in22;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_iftrue := VAR_in23;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_iffalse := VAR_in24;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_iftrue := VAR_in25;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iffalse := VAR_in26;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iftrue := VAR_in27;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iffalse := VAR_in28;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iftrue := VAR_in29;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iftrue := VAR_in3;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_iffalse := VAR_in30;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_iftrue := VAR_in31;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_iffalse := VAR_in32;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_iftrue := VAR_in33;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_iffalse := VAR_in34;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_iftrue := VAR_in35;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_iffalse := VAR_in36;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_iftrue := VAR_in37;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_iffalse := VAR_in38;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_iftrue := VAR_in39;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_iffalse := VAR_in4;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_iffalse := VAR_in40;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_iftrue := VAR_in41;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_iffalse := VAR_in42;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_iftrue := VAR_in43;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iffalse := VAR_in44;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iftrue := VAR_in45;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_iffalse := VAR_in46;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_iftrue := VAR_in47;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_iffalse := VAR_in48;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_iftrue := VAR_in49;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_iftrue := VAR_in5;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_iffalse := VAR_in50;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_iftrue := VAR_in51;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_iffalse := VAR_in52;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_iftrue := VAR_in53;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_iffalse := VAR_in54;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_iftrue := VAR_in55;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_iffalse := VAR_in56;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_iftrue := VAR_in57;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_iffalse := VAR_in58;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_iftrue := VAR_in59;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_iffalse := VAR_in6;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iffalse := VAR_in60;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iftrue := VAR_in61;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_iffalse := VAR_in62;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_iftrue := VAR_in63;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iffalse := VAR_in64;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iftrue := VAR_in65;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_iffalse := VAR_in66;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_iftrue := VAR_in67;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_iffalse := VAR_in68;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_iftrue := VAR_in69;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_iftrue := VAR_in7;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_iffalse := VAR_in70;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_iftrue := VAR_in71;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_iffalse := VAR_in72;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_iftrue := VAR_in73;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_iffalse := VAR_in74;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_iftrue := VAR_in75;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_iffalse := VAR_in76;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_iftrue := VAR_in77;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iffalse := VAR_in78;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iftrue := VAR_in79;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_iffalse := VAR_in8;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_iffalse := VAR_in80;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_iftrue := VAR_in81;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_iffalse := VAR_in82;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_iftrue := VAR_in83;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_iffalse := VAR_in84;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_iftrue := VAR_in85;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_iffalse := VAR_in86;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_iftrue := VAR_in87;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_iffalse := VAR_in88;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_iftrue := VAR_in89;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_iftrue := VAR_in9;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_iffalse := VAR_in90;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_iftrue := VAR_in91;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iffalse := VAR_in92;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iftrue := VAR_in93;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_iffalse := VAR_in94;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_iftrue := VAR_in95;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_iffalse := VAR_in96;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_iftrue := VAR_in97;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iffalse := VAR_in98;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iftrue := VAR_in99;
     -- uint7_2_2[bit_math_h_l1082_c10_1f09] LATENCY=0
     VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output := uint7_2_2(
     VAR_sel);

     -- uint7_4_4[bit_math_h_l1358_c10_c24c] LATENCY=0
     VAR_uint7_4_4_bit_math_h_l1358_c10_c24c_return_output := uint7_4_4(
     VAR_sel);

     -- uint7_3_3[bit_math_h_l1264_c10_78dc] LATENCY=0
     VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output := uint7_3_3(
     VAR_sel);

     -- uint7_5_5[bit_math_h_l1408_c10_901f] LATENCY=0
     VAR_uint7_5_5_bit_math_h_l1408_c10_901f_return_output := uint7_5_5(
     VAR_sel);

     -- uint7_6_6[bit_math_h_l1436_c10_87f9] LATENCY=0
     VAR_uint7_6_6_bit_math_h_l1436_c10_87f9_return_output := uint7_6_6(
     VAR_sel);

     -- uint7_1_1[bit_math_h_l724_c10_e4e1] LATENCY=0
     VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output := uint7_1_1(
     VAR_sel);

     -- uint7_0_0[bit_math_h_l14_c10_1a96] LATENCY=0
     VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output := uint7_0_0(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_cond := VAR_uint7_0_0_bit_math_h_l14_c10_1a96_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_cond := VAR_uint7_1_1_bit_math_h_l724_c10_e4e1_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_1f09_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_78dc_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_c24c_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_c24c_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_c24c_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_c24c_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_901f_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_901f_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_cond := VAR_uint7_6_6_bit_math_h_l1436_c10_87f9_return_output;
     -- layer0_node62_MUX[bit_math_h_l700_c3_0d13] LATENCY=0
     -- Inputs
     layer0_node62_MUX_bit_math_h_l700_c3_0d13_cond <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_cond;
     layer0_node62_MUX_bit_math_h_l700_c3_0d13_iftrue <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_iftrue;
     layer0_node62_MUX_bit_math_h_l700_c3_0d13_iffalse <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_iffalse;
     -- Outputs
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_return_output := layer0_node62_MUX_bit_math_h_l700_c3_0d13_return_output;

     -- layer0_node24_MUX[bit_math_h_l282_c3_670b] LATENCY=0
     -- Inputs
     layer0_node24_MUX_bit_math_h_l282_c3_670b_cond <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_cond;
     layer0_node24_MUX_bit_math_h_l282_c3_670b_iftrue <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_iftrue;
     layer0_node24_MUX_bit_math_h_l282_c3_670b_iffalse <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_iffalse;
     -- Outputs
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_return_output := layer0_node24_MUX_bit_math_h_l282_c3_670b_return_output;

     -- layer0_node53_MUX[bit_math_h_l601_c3_76ac] LATENCY=0
     -- Inputs
     layer0_node53_MUX_bit_math_h_l601_c3_76ac_cond <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_cond;
     layer0_node53_MUX_bit_math_h_l601_c3_76ac_iftrue <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_iftrue;
     layer0_node53_MUX_bit_math_h_l601_c3_76ac_iffalse <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_iffalse;
     -- Outputs
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_return_output := layer0_node53_MUX_bit_math_h_l601_c3_76ac_return_output;

     -- layer0_node55_MUX[bit_math_h_l623_c3_ec7e] LATENCY=0
     -- Inputs
     layer0_node55_MUX_bit_math_h_l623_c3_ec7e_cond <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_cond;
     layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iftrue <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iftrue;
     layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iffalse <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_iffalse;
     -- Outputs
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_return_output := layer0_node55_MUX_bit_math_h_l623_c3_ec7e_return_output;

     -- layer0_node29_MUX[bit_math_h_l337_c3_7a23] LATENCY=0
     -- Inputs
     layer0_node29_MUX_bit_math_h_l337_c3_7a23_cond <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_cond;
     layer0_node29_MUX_bit_math_h_l337_c3_7a23_iftrue <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_iftrue;
     layer0_node29_MUX_bit_math_h_l337_c3_7a23_iffalse <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_iffalse;
     -- Outputs
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_return_output := layer0_node29_MUX_bit_math_h_l337_c3_7a23_return_output;

     -- layer0_node5_MUX[bit_math_h_l73_c3_936b] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_936b_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_936b_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_936b_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_return_output := layer0_node5_MUX_bit_math_h_l73_c3_936b_return_output;

     -- layer0_node13_MUX[bit_math_h_l161_c3_3a1c] LATENCY=0
     -- Inputs
     layer0_node13_MUX_bit_math_h_l161_c3_3a1c_cond <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_cond;
     layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iftrue <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iftrue;
     layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iffalse <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_iffalse;
     -- Outputs
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_return_output := layer0_node13_MUX_bit_math_h_l161_c3_3a1c_return_output;

     -- layer0_node31_MUX[bit_math_h_l359_c3_208c] LATENCY=0
     -- Inputs
     layer0_node31_MUX_bit_math_h_l359_c3_208c_cond <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_cond;
     layer0_node31_MUX_bit_math_h_l359_c3_208c_iftrue <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_iftrue;
     layer0_node31_MUX_bit_math_h_l359_c3_208c_iffalse <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_iffalse;
     -- Outputs
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_return_output := layer0_node31_MUX_bit_math_h_l359_c3_208c_return_output;

     -- layer0_node49_MUX[bit_math_h_l557_c3_3c6d] LATENCY=0
     -- Inputs
     layer0_node49_MUX_bit_math_h_l557_c3_3c6d_cond <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_cond;
     layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iftrue <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iftrue;
     layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iffalse <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_iffalse;
     -- Outputs
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_return_output := layer0_node49_MUX_bit_math_h_l557_c3_3c6d_return_output;

     -- layer0_node61_MUX[bit_math_h_l689_c3_9f98] LATENCY=0
     -- Inputs
     layer0_node61_MUX_bit_math_h_l689_c3_9f98_cond <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_cond;
     layer0_node61_MUX_bit_math_h_l689_c3_9f98_iftrue <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_iftrue;
     layer0_node61_MUX_bit_math_h_l689_c3_9f98_iffalse <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_iffalse;
     -- Outputs
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_return_output := layer0_node61_MUX_bit_math_h_l689_c3_9f98_return_output;

     -- layer0_node18_MUX[bit_math_h_l216_c3_23c8] LATENCY=0
     -- Inputs
     layer0_node18_MUX_bit_math_h_l216_c3_23c8_cond <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_cond;
     layer0_node18_MUX_bit_math_h_l216_c3_23c8_iftrue <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_iftrue;
     layer0_node18_MUX_bit_math_h_l216_c3_23c8_iffalse <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_iffalse;
     -- Outputs
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_return_output := layer0_node18_MUX_bit_math_h_l216_c3_23c8_return_output;

     -- layer0_node47_MUX[bit_math_h_l535_c3_167a] LATENCY=0
     -- Inputs
     layer0_node47_MUX_bit_math_h_l535_c3_167a_cond <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_cond;
     layer0_node47_MUX_bit_math_h_l535_c3_167a_iftrue <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_iftrue;
     layer0_node47_MUX_bit_math_h_l535_c3_167a_iffalse <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_iffalse;
     -- Outputs
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_return_output := layer0_node47_MUX_bit_math_h_l535_c3_167a_return_output;

     -- layer0_node23_MUX[bit_math_h_l271_c3_6340] LATENCY=0
     -- Inputs
     layer0_node23_MUX_bit_math_h_l271_c3_6340_cond <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_cond;
     layer0_node23_MUX_bit_math_h_l271_c3_6340_iftrue <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_iftrue;
     layer0_node23_MUX_bit_math_h_l271_c3_6340_iffalse <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_iffalse;
     -- Outputs
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_return_output := layer0_node23_MUX_bit_math_h_l271_c3_6340_return_output;

     -- layer0_node51_MUX[bit_math_h_l579_c3_1b2f] LATENCY=0
     -- Inputs
     layer0_node51_MUX_bit_math_h_l579_c3_1b2f_cond <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_cond;
     layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iftrue <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iftrue;
     layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iffalse <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_iffalse;
     -- Outputs
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_return_output := layer0_node51_MUX_bit_math_h_l579_c3_1b2f_return_output;

     -- layer0_node60_MUX[bit_math_h_l678_c3_fe9f] LATENCY=0
     -- Inputs
     layer0_node60_MUX_bit_math_h_l678_c3_fe9f_cond <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_cond;
     layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iftrue <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iftrue;
     layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iffalse <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_iffalse;
     -- Outputs
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_return_output := layer0_node60_MUX_bit_math_h_l678_c3_fe9f_return_output;

     -- layer0_node1_MUX[bit_math_h_l29_c3_b2fc] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_b2fc_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_return_output := layer0_node1_MUX_bit_math_h_l29_c3_b2fc_return_output;

     -- layer0_node17_MUX[bit_math_h_l205_c3_39fd] LATENCY=0
     -- Inputs
     layer0_node17_MUX_bit_math_h_l205_c3_39fd_cond <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_cond;
     layer0_node17_MUX_bit_math_h_l205_c3_39fd_iftrue <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_iftrue;
     layer0_node17_MUX_bit_math_h_l205_c3_39fd_iffalse <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_iffalse;
     -- Outputs
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_return_output := layer0_node17_MUX_bit_math_h_l205_c3_39fd_return_output;

     -- layer0_node63_MUX[bit_math_h_l711_c3_2778] LATENCY=0
     -- Inputs
     layer0_node63_MUX_bit_math_h_l711_c3_2778_cond <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_cond;
     layer0_node63_MUX_bit_math_h_l711_c3_2778_iftrue <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_iftrue;
     layer0_node63_MUX_bit_math_h_l711_c3_2778_iffalse <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_iffalse;
     -- Outputs
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_return_output := layer0_node63_MUX_bit_math_h_l711_c3_2778_return_output;

     -- layer0_node10_MUX[bit_math_h_l128_c3_0e40] LATENCY=0
     -- Inputs
     layer0_node10_MUX_bit_math_h_l128_c3_0e40_cond <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_cond;
     layer0_node10_MUX_bit_math_h_l128_c3_0e40_iftrue <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_iftrue;
     layer0_node10_MUX_bit_math_h_l128_c3_0e40_iffalse <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_iffalse;
     -- Outputs
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_return_output := layer0_node10_MUX_bit_math_h_l128_c3_0e40_return_output;

     -- layer0_node43_MUX[bit_math_h_l491_c3_001b] LATENCY=0
     -- Inputs
     layer0_node43_MUX_bit_math_h_l491_c3_001b_cond <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_cond;
     layer0_node43_MUX_bit_math_h_l491_c3_001b_iftrue <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_iftrue;
     layer0_node43_MUX_bit_math_h_l491_c3_001b_iffalse <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_iffalse;
     -- Outputs
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_return_output := layer0_node43_MUX_bit_math_h_l491_c3_001b_return_output;

     -- layer0_node27_MUX[bit_math_h_l315_c3_ac24] LATENCY=0
     -- Inputs
     layer0_node27_MUX_bit_math_h_l315_c3_ac24_cond <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_cond;
     layer0_node27_MUX_bit_math_h_l315_c3_ac24_iftrue <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_iftrue;
     layer0_node27_MUX_bit_math_h_l315_c3_ac24_iffalse <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_iffalse;
     -- Outputs
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_return_output := layer0_node27_MUX_bit_math_h_l315_c3_ac24_return_output;

     -- layer0_node39_MUX[bit_math_h_l447_c3_b0c4] LATENCY=0
     -- Inputs
     layer0_node39_MUX_bit_math_h_l447_c3_b0c4_cond <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_cond;
     layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iftrue <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iftrue;
     layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iffalse <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_iffalse;
     -- Outputs
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_return_output := layer0_node39_MUX_bit_math_h_l447_c3_b0c4_return_output;

     -- layer0_node54_MUX[bit_math_h_l612_c3_e1c8] LATENCY=0
     -- Inputs
     layer0_node54_MUX_bit_math_h_l612_c3_e1c8_cond <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_cond;
     layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iftrue <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iftrue;
     layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iffalse <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_iffalse;
     -- Outputs
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_return_output := layer0_node54_MUX_bit_math_h_l612_c3_e1c8_return_output;

     -- layer0_node19_MUX[bit_math_h_l227_c3_ea58] LATENCY=0
     -- Inputs
     layer0_node19_MUX_bit_math_h_l227_c3_ea58_cond <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_cond;
     layer0_node19_MUX_bit_math_h_l227_c3_ea58_iftrue <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_iftrue;
     layer0_node19_MUX_bit_math_h_l227_c3_ea58_iffalse <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_iffalse;
     -- Outputs
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_return_output := layer0_node19_MUX_bit_math_h_l227_c3_ea58_return_output;

     -- layer0_node36_MUX[bit_math_h_l414_c3_0db7] LATENCY=0
     -- Inputs
     layer0_node36_MUX_bit_math_h_l414_c3_0db7_cond <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_cond;
     layer0_node36_MUX_bit_math_h_l414_c3_0db7_iftrue <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_iftrue;
     layer0_node36_MUX_bit_math_h_l414_c3_0db7_iffalse <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_iffalse;
     -- Outputs
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_return_output := layer0_node36_MUX_bit_math_h_l414_c3_0db7_return_output;

     -- layer0_node35_MUX[bit_math_h_l403_c3_749b] LATENCY=0
     -- Inputs
     layer0_node35_MUX_bit_math_h_l403_c3_749b_cond <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_cond;
     layer0_node35_MUX_bit_math_h_l403_c3_749b_iftrue <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_iftrue;
     layer0_node35_MUX_bit_math_h_l403_c3_749b_iffalse <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_iffalse;
     -- Outputs
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_return_output := layer0_node35_MUX_bit_math_h_l403_c3_749b_return_output;

     -- layer0_node37_MUX[bit_math_h_l425_c3_7f65] LATENCY=0
     -- Inputs
     layer0_node37_MUX_bit_math_h_l425_c3_7f65_cond <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_cond;
     layer0_node37_MUX_bit_math_h_l425_c3_7f65_iftrue <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_iftrue;
     layer0_node37_MUX_bit_math_h_l425_c3_7f65_iffalse <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_iffalse;
     -- Outputs
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_return_output := layer0_node37_MUX_bit_math_h_l425_c3_7f65_return_output;

     -- layer0_node41_MUX[bit_math_h_l469_c3_62cc] LATENCY=0
     -- Inputs
     layer0_node41_MUX_bit_math_h_l469_c3_62cc_cond <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_cond;
     layer0_node41_MUX_bit_math_h_l469_c3_62cc_iftrue <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_iftrue;
     layer0_node41_MUX_bit_math_h_l469_c3_62cc_iffalse <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_iffalse;
     -- Outputs
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_return_output := layer0_node41_MUX_bit_math_h_l469_c3_62cc_return_output;

     -- layer0_node33_MUX[bit_math_h_l381_c3_0aac] LATENCY=0
     -- Inputs
     layer0_node33_MUX_bit_math_h_l381_c3_0aac_cond <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_cond;
     layer0_node33_MUX_bit_math_h_l381_c3_0aac_iftrue <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_iftrue;
     layer0_node33_MUX_bit_math_h_l381_c3_0aac_iffalse <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_iffalse;
     -- Outputs
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_return_output := layer0_node33_MUX_bit_math_h_l381_c3_0aac_return_output;

     -- layer0_node40_MUX[bit_math_h_l458_c3_773e] LATENCY=0
     -- Inputs
     layer0_node40_MUX_bit_math_h_l458_c3_773e_cond <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_cond;
     layer0_node40_MUX_bit_math_h_l458_c3_773e_iftrue <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_iftrue;
     layer0_node40_MUX_bit_math_h_l458_c3_773e_iffalse <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_iffalse;
     -- Outputs
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_return_output := layer0_node40_MUX_bit_math_h_l458_c3_773e_return_output;

     -- layer0_node15_MUX[bit_math_h_l183_c3_392b] LATENCY=0
     -- Inputs
     layer0_node15_MUX_bit_math_h_l183_c3_392b_cond <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_cond;
     layer0_node15_MUX_bit_math_h_l183_c3_392b_iftrue <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_iftrue;
     layer0_node15_MUX_bit_math_h_l183_c3_392b_iffalse <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_iffalse;
     -- Outputs
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_return_output := layer0_node15_MUX_bit_math_h_l183_c3_392b_return_output;

     -- layer0_node14_MUX[bit_math_h_l172_c3_7ef7] LATENCY=0
     -- Inputs
     layer0_node14_MUX_bit_math_h_l172_c3_7ef7_cond <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_cond;
     layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iftrue <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iftrue;
     layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iffalse <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_iffalse;
     -- Outputs
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_return_output := layer0_node14_MUX_bit_math_h_l172_c3_7ef7_return_output;

     -- layer0_node12_MUX[bit_math_h_l150_c3_1560] LATENCY=0
     -- Inputs
     layer0_node12_MUX_bit_math_h_l150_c3_1560_cond <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_cond;
     layer0_node12_MUX_bit_math_h_l150_c3_1560_iftrue <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_iftrue;
     layer0_node12_MUX_bit_math_h_l150_c3_1560_iffalse <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_iffalse;
     -- Outputs
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_return_output := layer0_node12_MUX_bit_math_h_l150_c3_1560_return_output;

     -- layer0_node22_MUX[bit_math_h_l260_c3_1c3c] LATENCY=0
     -- Inputs
     layer0_node22_MUX_bit_math_h_l260_c3_1c3c_cond <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_cond;
     layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iftrue <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iftrue;
     layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iffalse <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_iffalse;
     -- Outputs
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_return_output := layer0_node22_MUX_bit_math_h_l260_c3_1c3c_return_output;

     -- layer0_node58_MUX[bit_math_h_l656_c3_e8c0] LATENCY=0
     -- Inputs
     layer0_node58_MUX_bit_math_h_l656_c3_e8c0_cond <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_cond;
     layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iftrue <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iftrue;
     layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iffalse <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_iffalse;
     -- Outputs
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_return_output := layer0_node58_MUX_bit_math_h_l656_c3_e8c0_return_output;

     -- layer0_node57_MUX[bit_math_h_l645_c3_d7f5] LATENCY=0
     -- Inputs
     layer0_node57_MUX_bit_math_h_l645_c3_d7f5_cond <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_cond;
     layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iftrue <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iftrue;
     layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iffalse <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_iffalse;
     -- Outputs
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_return_output := layer0_node57_MUX_bit_math_h_l645_c3_d7f5_return_output;

     -- layer0_node20_MUX[bit_math_h_l238_c3_eb78] LATENCY=0
     -- Inputs
     layer0_node20_MUX_bit_math_h_l238_c3_eb78_cond <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_cond;
     layer0_node20_MUX_bit_math_h_l238_c3_eb78_iftrue <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_iftrue;
     layer0_node20_MUX_bit_math_h_l238_c3_eb78_iffalse <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_iffalse;
     -- Outputs
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_return_output := layer0_node20_MUX_bit_math_h_l238_c3_eb78_return_output;

     -- layer0_node32_MUX[bit_math_h_l370_c3_bcd8] LATENCY=0
     -- Inputs
     layer0_node32_MUX_bit_math_h_l370_c3_bcd8_cond <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_cond;
     layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iftrue <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iftrue;
     layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iffalse <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_iffalse;
     -- Outputs
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_return_output := layer0_node32_MUX_bit_math_h_l370_c3_bcd8_return_output;

     -- layer0_node42_MUX[bit_math_h_l480_c3_d626] LATENCY=0
     -- Inputs
     layer0_node42_MUX_bit_math_h_l480_c3_d626_cond <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_cond;
     layer0_node42_MUX_bit_math_h_l480_c3_d626_iftrue <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_iftrue;
     layer0_node42_MUX_bit_math_h_l480_c3_d626_iffalse <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_iffalse;
     -- Outputs
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_return_output := layer0_node42_MUX_bit_math_h_l480_c3_d626_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_f259] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_f259_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_f259_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_f259_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_return_output := layer0_node7_MUX_bit_math_h_l95_c3_f259_return_output;

     -- layer0_node30_MUX[bit_math_h_l348_c3_7ed3] LATENCY=0
     -- Inputs
     layer0_node30_MUX_bit_math_h_l348_c3_7ed3_cond <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_cond;
     layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iftrue <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iftrue;
     layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iffalse <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_iffalse;
     -- Outputs
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_return_output := layer0_node30_MUX_bit_math_h_l348_c3_7ed3_return_output;

     -- layer0_node50_MUX[bit_math_h_l568_c3_e0e2] LATENCY=0
     -- Inputs
     layer0_node50_MUX_bit_math_h_l568_c3_e0e2_cond <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_cond;
     layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iftrue <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iftrue;
     layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iffalse <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_iffalse;
     -- Outputs
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_return_output := layer0_node50_MUX_bit_math_h_l568_c3_e0e2_return_output;

     -- layer0_node45_MUX[bit_math_h_l513_c3_cc83] LATENCY=0
     -- Inputs
     layer0_node45_MUX_bit_math_h_l513_c3_cc83_cond <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_cond;
     layer0_node45_MUX_bit_math_h_l513_c3_cc83_iftrue <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_iftrue;
     layer0_node45_MUX_bit_math_h_l513_c3_cc83_iffalse <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_iffalse;
     -- Outputs
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_return_output := layer0_node45_MUX_bit_math_h_l513_c3_cc83_return_output;

     -- layer0_node11_MUX[bit_math_h_l139_c3_381c] LATENCY=0
     -- Inputs
     layer0_node11_MUX_bit_math_h_l139_c3_381c_cond <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_cond;
     layer0_node11_MUX_bit_math_h_l139_c3_381c_iftrue <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_iftrue;
     layer0_node11_MUX_bit_math_h_l139_c3_381c_iffalse <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_iffalse;
     -- Outputs
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_return_output := layer0_node11_MUX_bit_math_h_l139_c3_381c_return_output;

     -- layer0_node6_MUX[bit_math_h_l84_c3_6f9a] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_6f9a_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_return_output := layer0_node6_MUX_bit_math_h_l84_c3_6f9a_return_output;

     -- layer0_node16_MUX[bit_math_h_l194_c3_cada] LATENCY=0
     -- Inputs
     layer0_node16_MUX_bit_math_h_l194_c3_cada_cond <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_cond;
     layer0_node16_MUX_bit_math_h_l194_c3_cada_iftrue <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_iftrue;
     layer0_node16_MUX_bit_math_h_l194_c3_cada_iffalse <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_iffalse;
     -- Outputs
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_return_output := layer0_node16_MUX_bit_math_h_l194_c3_cada_return_output;

     -- layer0_node38_MUX[bit_math_h_l436_c3_d774] LATENCY=0
     -- Inputs
     layer0_node38_MUX_bit_math_h_l436_c3_d774_cond <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_cond;
     layer0_node38_MUX_bit_math_h_l436_c3_d774_iftrue <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_iftrue;
     layer0_node38_MUX_bit_math_h_l436_c3_d774_iffalse <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_iffalse;
     -- Outputs
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_return_output := layer0_node38_MUX_bit_math_h_l436_c3_d774_return_output;

     -- layer0_node26_MUX[bit_math_h_l304_c3_53e2] LATENCY=0
     -- Inputs
     layer0_node26_MUX_bit_math_h_l304_c3_53e2_cond <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_cond;
     layer0_node26_MUX_bit_math_h_l304_c3_53e2_iftrue <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_iftrue;
     layer0_node26_MUX_bit_math_h_l304_c3_53e2_iffalse <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_iffalse;
     -- Outputs
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_return_output := layer0_node26_MUX_bit_math_h_l304_c3_53e2_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_be4c] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_be4c_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_be4c_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_be4c_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_return_output := layer0_node4_MUX_bit_math_h_l62_c3_be4c_return_output;

     -- layer0_node28_MUX[bit_math_h_l326_c3_97ed] LATENCY=0
     -- Inputs
     layer0_node28_MUX_bit_math_h_l326_c3_97ed_cond <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_cond;
     layer0_node28_MUX_bit_math_h_l326_c3_97ed_iftrue <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_iftrue;
     layer0_node28_MUX_bit_math_h_l326_c3_97ed_iffalse <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_iffalse;
     -- Outputs
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_return_output := layer0_node28_MUX_bit_math_h_l326_c3_97ed_return_output;

     -- layer0_node9_MUX[bit_math_h_l117_c3_1a47] LATENCY=0
     -- Inputs
     layer0_node9_MUX_bit_math_h_l117_c3_1a47_cond <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_cond;
     layer0_node9_MUX_bit_math_h_l117_c3_1a47_iftrue <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_iftrue;
     layer0_node9_MUX_bit_math_h_l117_c3_1a47_iffalse <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_iffalse;
     -- Outputs
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_return_output := layer0_node9_MUX_bit_math_h_l117_c3_1a47_return_output;

     -- layer0_node48_MUX[bit_math_h_l546_c3_41a2] LATENCY=0
     -- Inputs
     layer0_node48_MUX_bit_math_h_l546_c3_41a2_cond <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_cond;
     layer0_node48_MUX_bit_math_h_l546_c3_41a2_iftrue <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_iftrue;
     layer0_node48_MUX_bit_math_h_l546_c3_41a2_iffalse <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_iffalse;
     -- Outputs
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_return_output := layer0_node48_MUX_bit_math_h_l546_c3_41a2_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_13b9] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_13b9_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_13b9_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_13b9_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_return_output := layer0_node3_MUX_bit_math_h_l51_c3_13b9_return_output;

     -- layer0_node44_MUX[bit_math_h_l502_c3_1816] LATENCY=0
     -- Inputs
     layer0_node44_MUX_bit_math_h_l502_c3_1816_cond <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_cond;
     layer0_node44_MUX_bit_math_h_l502_c3_1816_iftrue <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_iftrue;
     layer0_node44_MUX_bit_math_h_l502_c3_1816_iffalse <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_iffalse;
     -- Outputs
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_return_output := layer0_node44_MUX_bit_math_h_l502_c3_1816_return_output;

     -- layer0_node21_MUX[bit_math_h_l249_c3_228d] LATENCY=0
     -- Inputs
     layer0_node21_MUX_bit_math_h_l249_c3_228d_cond <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_cond;
     layer0_node21_MUX_bit_math_h_l249_c3_228d_iftrue <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_iftrue;
     layer0_node21_MUX_bit_math_h_l249_c3_228d_iffalse <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_iffalse;
     -- Outputs
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_return_output := layer0_node21_MUX_bit_math_h_l249_c3_228d_return_output;

     -- layer0_node52_MUX[bit_math_h_l590_c3_dee1] LATENCY=0
     -- Inputs
     layer0_node52_MUX_bit_math_h_l590_c3_dee1_cond <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_cond;
     layer0_node52_MUX_bit_math_h_l590_c3_dee1_iftrue <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_iftrue;
     layer0_node52_MUX_bit_math_h_l590_c3_dee1_iffalse <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_iffalse;
     -- Outputs
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_return_output := layer0_node52_MUX_bit_math_h_l590_c3_dee1_return_output;

     -- layer0_node46_MUX[bit_math_h_l524_c3_aa0a] LATENCY=0
     -- Inputs
     layer0_node46_MUX_bit_math_h_l524_c3_aa0a_cond <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_cond;
     layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iftrue <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iftrue;
     layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iffalse <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_iffalse;
     -- Outputs
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_return_output := layer0_node46_MUX_bit_math_h_l524_c3_aa0a_return_output;

     -- layer0_node34_MUX[bit_math_h_l392_c3_6801] LATENCY=0
     -- Inputs
     layer0_node34_MUX_bit_math_h_l392_c3_6801_cond <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_cond;
     layer0_node34_MUX_bit_math_h_l392_c3_6801_iftrue <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_iftrue;
     layer0_node34_MUX_bit_math_h_l392_c3_6801_iffalse <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_iffalse;
     -- Outputs
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_return_output := layer0_node34_MUX_bit_math_h_l392_c3_6801_return_output;

     -- layer0_node25_MUX[bit_math_h_l293_c3_83e8] LATENCY=0
     -- Inputs
     layer0_node25_MUX_bit_math_h_l293_c3_83e8_cond <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_cond;
     layer0_node25_MUX_bit_math_h_l293_c3_83e8_iftrue <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_iftrue;
     layer0_node25_MUX_bit_math_h_l293_c3_83e8_iffalse <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_iffalse;
     -- Outputs
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_return_output := layer0_node25_MUX_bit_math_h_l293_c3_83e8_return_output;

     -- layer0_node59_MUX[bit_math_h_l667_c3_1ea2] LATENCY=0
     -- Inputs
     layer0_node59_MUX_bit_math_h_l667_c3_1ea2_cond <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_cond;
     layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iftrue <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iftrue;
     layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iffalse <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_iffalse;
     -- Outputs
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_return_output := layer0_node59_MUX_bit_math_h_l667_c3_1ea2_return_output;

     -- layer0_node8_MUX[bit_math_h_l106_c3_2e0c] LATENCY=0
     -- Inputs
     layer0_node8_MUX_bit_math_h_l106_c3_2e0c_cond <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_cond;
     layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iftrue <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iftrue;
     layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iffalse <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_iffalse;
     -- Outputs
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_return_output := layer0_node8_MUX_bit_math_h_l106_c3_2e0c_return_output;

     -- layer0_node56_MUX[bit_math_h_l634_c3_5b10] LATENCY=0
     -- Inputs
     layer0_node56_MUX_bit_math_h_l634_c3_5b10_cond <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_cond;
     layer0_node56_MUX_bit_math_h_l634_c3_5b10_iftrue <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_iftrue;
     layer0_node56_MUX_bit_math_h_l634_c3_5b10_iffalse <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_iffalse;
     -- Outputs
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_return_output := layer0_node56_MUX_bit_math_h_l634_c3_5b10_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_3d12] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_3d12_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_3d12_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_3d12_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_return_output := layer0_node2_MUX_bit_math_h_l40_c3_3d12_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_8bd4] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_8bd4_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_return_output := layer0_node0_MUX_bit_math_h_l18_c3_8bd4_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_8bd4_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_iffalse := VAR_layer0_node10_MUX_bit_math_h_l128_c3_0e40_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_iftrue := VAR_layer0_node11_MUX_bit_math_h_l139_c3_381c_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_iffalse := VAR_layer0_node12_MUX_bit_math_h_l150_c3_1560_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_iftrue := VAR_layer0_node13_MUX_bit_math_h_l161_c3_3a1c_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iffalse := VAR_layer0_node14_MUX_bit_math_h_l172_c3_7ef7_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iftrue := VAR_layer0_node15_MUX_bit_math_h_l183_c3_392b_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_iffalse := VAR_layer0_node16_MUX_bit_math_h_l194_c3_cada_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_iftrue := VAR_layer0_node17_MUX_bit_math_h_l205_c3_39fd_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_iffalse := VAR_layer0_node18_MUX_bit_math_h_l216_c3_23c8_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_iftrue := VAR_layer0_node19_MUX_bit_math_h_l227_c3_ea58_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_b2fc_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_iffalse := VAR_layer0_node20_MUX_bit_math_h_l238_c3_eb78_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_iftrue := VAR_layer0_node21_MUX_bit_math_h_l249_c3_228d_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_iffalse := VAR_layer0_node22_MUX_bit_math_h_l260_c3_1c3c_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_iftrue := VAR_layer0_node23_MUX_bit_math_h_l271_c3_6340_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_iffalse := VAR_layer0_node24_MUX_bit_math_h_l282_c3_670b_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_iftrue := VAR_layer0_node25_MUX_bit_math_h_l293_c3_83e8_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iffalse := VAR_layer0_node26_MUX_bit_math_h_l304_c3_53e2_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iftrue := VAR_layer0_node27_MUX_bit_math_h_l315_c3_ac24_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_iffalse := VAR_layer0_node28_MUX_bit_math_h_l326_c3_97ed_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_iftrue := VAR_layer0_node29_MUX_bit_math_h_l337_c3_7a23_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_3d12_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_iffalse := VAR_layer0_node30_MUX_bit_math_h_l348_c3_7ed3_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_iftrue := VAR_layer0_node31_MUX_bit_math_h_l359_c3_208c_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iffalse := VAR_layer0_node32_MUX_bit_math_h_l370_c3_bcd8_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iftrue := VAR_layer0_node33_MUX_bit_math_h_l381_c3_0aac_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_iffalse := VAR_layer0_node34_MUX_bit_math_h_l392_c3_6801_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_iftrue := VAR_layer0_node35_MUX_bit_math_h_l403_c3_749b_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iffalse := VAR_layer0_node36_MUX_bit_math_h_l414_c3_0db7_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iftrue := VAR_layer0_node37_MUX_bit_math_h_l425_c3_7f65_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_iffalse := VAR_layer0_node38_MUX_bit_math_h_l436_c3_d774_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_iftrue := VAR_layer0_node39_MUX_bit_math_h_l447_c3_b0c4_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_13b9_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iffalse := VAR_layer0_node40_MUX_bit_math_h_l458_c3_773e_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iftrue := VAR_layer0_node41_MUX_bit_math_h_l469_c3_62cc_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_iffalse := VAR_layer0_node42_MUX_bit_math_h_l480_c3_d626_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_iftrue := VAR_layer0_node43_MUX_bit_math_h_l491_c3_001b_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iffalse := VAR_layer0_node44_MUX_bit_math_h_l502_c3_1816_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iftrue := VAR_layer0_node45_MUX_bit_math_h_l513_c3_cc83_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iffalse := VAR_layer0_node46_MUX_bit_math_h_l524_c3_aa0a_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iftrue := VAR_layer0_node47_MUX_bit_math_h_l535_c3_167a_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_iffalse := VAR_layer0_node48_MUX_bit_math_h_l546_c3_41a2_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_iftrue := VAR_layer0_node49_MUX_bit_math_h_l557_c3_3c6d_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_be4c_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iffalse := VAR_layer0_node50_MUX_bit_math_h_l568_c3_e0e2_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iftrue := VAR_layer0_node51_MUX_bit_math_h_l579_c3_1b2f_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iffalse := VAR_layer0_node52_MUX_bit_math_h_l590_c3_dee1_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iftrue := VAR_layer0_node53_MUX_bit_math_h_l601_c3_76ac_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iffalse := VAR_layer0_node54_MUX_bit_math_h_l612_c3_e1c8_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iftrue := VAR_layer0_node55_MUX_bit_math_h_l623_c3_ec7e_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_iffalse := VAR_layer0_node56_MUX_bit_math_h_l634_c3_5b10_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_iftrue := VAR_layer0_node57_MUX_bit_math_h_l645_c3_d7f5_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iffalse := VAR_layer0_node58_MUX_bit_math_h_l656_c3_e8c0_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iftrue := VAR_layer0_node59_MUX_bit_math_h_l667_c3_1ea2_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_936b_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iffalse := VAR_layer0_node60_MUX_bit_math_h_l678_c3_fe9f_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iftrue := VAR_layer0_node61_MUX_bit_math_h_l689_c3_9f98_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iffalse := VAR_layer0_node62_MUX_bit_math_h_l700_c3_0d13_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iftrue := VAR_layer0_node63_MUX_bit_math_h_l711_c3_2778_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_6f9a_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_f259_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_iffalse := VAR_layer0_node8_MUX_bit_math_h_l106_c3_2e0c_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_iftrue := VAR_layer0_node9_MUX_bit_math_h_l117_c3_1a47_return_output;
     -- layer1_node23_MUX[bit_math_h_l981_c3_d2b9] LATENCY=0
     -- Inputs
     layer1_node23_MUX_bit_math_h_l981_c3_d2b9_cond <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_cond;
     layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iftrue <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iftrue;
     layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iffalse <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_iffalse;
     -- Outputs
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_return_output := layer1_node23_MUX_bit_math_h_l981_c3_d2b9_return_output;

     -- layer1_node14_MUX[bit_math_h_l882_c3_9be0] LATENCY=0
     -- Inputs
     layer1_node14_MUX_bit_math_h_l882_c3_9be0_cond <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_cond;
     layer1_node14_MUX_bit_math_h_l882_c3_9be0_iftrue <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_iftrue;
     layer1_node14_MUX_bit_math_h_l882_c3_9be0_iffalse <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_iffalse;
     -- Outputs
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_return_output := layer1_node14_MUX_bit_math_h_l882_c3_9be0_return_output;

     -- layer1_node1_MUX[bit_math_h_l739_c3_5e54] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l739_c3_5e54_cond <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_cond;
     layer1_node1_MUX_bit_math_h_l739_c3_5e54_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_iftrue;
     layer1_node1_MUX_bit_math_h_l739_c3_5e54_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_return_output := layer1_node1_MUX_bit_math_h_l739_c3_5e54_return_output;

     -- layer1_node13_MUX[bit_math_h_l871_c3_9f0e] LATENCY=0
     -- Inputs
     layer1_node13_MUX_bit_math_h_l871_c3_9f0e_cond <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_cond;
     layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iftrue <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iftrue;
     layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iffalse <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_iffalse;
     -- Outputs
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_return_output := layer1_node13_MUX_bit_math_h_l871_c3_9f0e_return_output;

     -- layer1_node11_MUX[bit_math_h_l849_c3_0669] LATENCY=0
     -- Inputs
     layer1_node11_MUX_bit_math_h_l849_c3_0669_cond <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_cond;
     layer1_node11_MUX_bit_math_h_l849_c3_0669_iftrue <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_iftrue;
     layer1_node11_MUX_bit_math_h_l849_c3_0669_iffalse <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_iffalse;
     -- Outputs
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_return_output := layer1_node11_MUX_bit_math_h_l849_c3_0669_return_output;

     -- layer1_node26_MUX[bit_math_h_l1014_c3_f8c1] LATENCY=0
     -- Inputs
     layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_cond <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_cond;
     layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iftrue <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iftrue;
     layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iffalse <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_iffalse;
     -- Outputs
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_return_output := layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_return_output;

     -- layer1_node24_MUX[bit_math_h_l992_c3_8792] LATENCY=0
     -- Inputs
     layer1_node24_MUX_bit_math_h_l992_c3_8792_cond <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_cond;
     layer1_node24_MUX_bit_math_h_l992_c3_8792_iftrue <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_iftrue;
     layer1_node24_MUX_bit_math_h_l992_c3_8792_iffalse <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_iffalse;
     -- Outputs
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_return_output := layer1_node24_MUX_bit_math_h_l992_c3_8792_return_output;

     -- layer1_node5_MUX[bit_math_h_l783_c3_7132] LATENCY=0
     -- Inputs
     layer1_node5_MUX_bit_math_h_l783_c3_7132_cond <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_cond;
     layer1_node5_MUX_bit_math_h_l783_c3_7132_iftrue <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_iftrue;
     layer1_node5_MUX_bit_math_h_l783_c3_7132_iffalse <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_iffalse;
     -- Outputs
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_return_output := layer1_node5_MUX_bit_math_h_l783_c3_7132_return_output;

     -- layer1_node4_MUX[bit_math_h_l772_c3_535b] LATENCY=0
     -- Inputs
     layer1_node4_MUX_bit_math_h_l772_c3_535b_cond <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_cond;
     layer1_node4_MUX_bit_math_h_l772_c3_535b_iftrue <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_iftrue;
     layer1_node4_MUX_bit_math_h_l772_c3_535b_iffalse <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_iffalse;
     -- Outputs
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_return_output := layer1_node4_MUX_bit_math_h_l772_c3_535b_return_output;

     -- layer1_node30_MUX[bit_math_h_l1058_c3_d1f5] LATENCY=0
     -- Inputs
     layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_cond <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_cond;
     layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iftrue <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iftrue;
     layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iffalse <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_iffalse;
     -- Outputs
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_return_output := layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_return_output;

     -- layer1_node28_MUX[bit_math_h_l1036_c3_deef] LATENCY=0
     -- Inputs
     layer1_node28_MUX_bit_math_h_l1036_c3_deef_cond <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_cond;
     layer1_node28_MUX_bit_math_h_l1036_c3_deef_iftrue <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_iftrue;
     layer1_node28_MUX_bit_math_h_l1036_c3_deef_iffalse <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_iffalse;
     -- Outputs
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_return_output := layer1_node28_MUX_bit_math_h_l1036_c3_deef_return_output;

     -- layer1_node2_MUX[bit_math_h_l750_c3_386d] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l750_c3_386d_cond <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_cond;
     layer1_node2_MUX_bit_math_h_l750_c3_386d_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_iftrue;
     layer1_node2_MUX_bit_math_h_l750_c3_386d_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_return_output := layer1_node2_MUX_bit_math_h_l750_c3_386d_return_output;

     -- layer1_node22_MUX[bit_math_h_l970_c3_3aa5] LATENCY=0
     -- Inputs
     layer1_node22_MUX_bit_math_h_l970_c3_3aa5_cond <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_cond;
     layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iftrue <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iftrue;
     layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iffalse <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_iffalse;
     -- Outputs
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_return_output := layer1_node22_MUX_bit_math_h_l970_c3_3aa5_return_output;

     -- layer1_node7_MUX[bit_math_h_l805_c3_a7b7] LATENCY=0
     -- Inputs
     layer1_node7_MUX_bit_math_h_l805_c3_a7b7_cond <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_cond;
     layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iftrue <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iftrue;
     layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iffalse <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_iffalse;
     -- Outputs
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_return_output := layer1_node7_MUX_bit_math_h_l805_c3_a7b7_return_output;

     -- layer1_node3_MUX[bit_math_h_l761_c3_c96d] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l761_c3_c96d_cond <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_cond;
     layer1_node3_MUX_bit_math_h_l761_c3_c96d_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_iftrue;
     layer1_node3_MUX_bit_math_h_l761_c3_c96d_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_return_output := layer1_node3_MUX_bit_math_h_l761_c3_c96d_return_output;

     -- layer1_node16_MUX[bit_math_h_l904_c3_fdb3] LATENCY=0
     -- Inputs
     layer1_node16_MUX_bit_math_h_l904_c3_fdb3_cond <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_cond;
     layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iftrue <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iftrue;
     layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iffalse <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_iffalse;
     -- Outputs
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_return_output := layer1_node16_MUX_bit_math_h_l904_c3_fdb3_return_output;

     -- layer1_node19_MUX[bit_math_h_l937_c3_1a24] LATENCY=0
     -- Inputs
     layer1_node19_MUX_bit_math_h_l937_c3_1a24_cond <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_cond;
     layer1_node19_MUX_bit_math_h_l937_c3_1a24_iftrue <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_iftrue;
     layer1_node19_MUX_bit_math_h_l937_c3_1a24_iffalse <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_iffalse;
     -- Outputs
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_return_output := layer1_node19_MUX_bit_math_h_l937_c3_1a24_return_output;

     -- layer1_node20_MUX[bit_math_h_l948_c3_2dbc] LATENCY=0
     -- Inputs
     layer1_node20_MUX_bit_math_h_l948_c3_2dbc_cond <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_cond;
     layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iftrue <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iftrue;
     layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iffalse <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_iffalse;
     -- Outputs
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_return_output := layer1_node20_MUX_bit_math_h_l948_c3_2dbc_return_output;

     -- layer1_node17_MUX[bit_math_h_l915_c3_bba5] LATENCY=0
     -- Inputs
     layer1_node17_MUX_bit_math_h_l915_c3_bba5_cond <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_cond;
     layer1_node17_MUX_bit_math_h_l915_c3_bba5_iftrue <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_iftrue;
     layer1_node17_MUX_bit_math_h_l915_c3_bba5_iffalse <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_iffalse;
     -- Outputs
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_return_output := layer1_node17_MUX_bit_math_h_l915_c3_bba5_return_output;

     -- layer1_node9_MUX[bit_math_h_l827_c3_90fc] LATENCY=0
     -- Inputs
     layer1_node9_MUX_bit_math_h_l827_c3_90fc_cond <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_cond;
     layer1_node9_MUX_bit_math_h_l827_c3_90fc_iftrue <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_iftrue;
     layer1_node9_MUX_bit_math_h_l827_c3_90fc_iffalse <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_iffalse;
     -- Outputs
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_return_output := layer1_node9_MUX_bit_math_h_l827_c3_90fc_return_output;

     -- layer1_node29_MUX[bit_math_h_l1047_c3_d4d6] LATENCY=0
     -- Inputs
     layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_cond <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_cond;
     layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iftrue <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iftrue;
     layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iffalse <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_iffalse;
     -- Outputs
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_return_output := layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_return_output;

     -- layer1_node25_MUX[bit_math_h_l1003_c3_2c90] LATENCY=0
     -- Inputs
     layer1_node25_MUX_bit_math_h_l1003_c3_2c90_cond <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_cond;
     layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iftrue <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iftrue;
     layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iffalse <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_iffalse;
     -- Outputs
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_return_output := layer1_node25_MUX_bit_math_h_l1003_c3_2c90_return_output;

     -- layer1_node21_MUX[bit_math_h_l959_c3_f718] LATENCY=0
     -- Inputs
     layer1_node21_MUX_bit_math_h_l959_c3_f718_cond <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_cond;
     layer1_node21_MUX_bit_math_h_l959_c3_f718_iftrue <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_iftrue;
     layer1_node21_MUX_bit_math_h_l959_c3_f718_iffalse <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_iffalse;
     -- Outputs
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_return_output := layer1_node21_MUX_bit_math_h_l959_c3_f718_return_output;

     -- layer1_node15_MUX[bit_math_h_l893_c3_db88] LATENCY=0
     -- Inputs
     layer1_node15_MUX_bit_math_h_l893_c3_db88_cond <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_cond;
     layer1_node15_MUX_bit_math_h_l893_c3_db88_iftrue <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_iftrue;
     layer1_node15_MUX_bit_math_h_l893_c3_db88_iffalse <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_iffalse;
     -- Outputs
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_return_output := layer1_node15_MUX_bit_math_h_l893_c3_db88_return_output;

     -- layer1_node12_MUX[bit_math_h_l860_c3_f017] LATENCY=0
     -- Inputs
     layer1_node12_MUX_bit_math_h_l860_c3_f017_cond <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_cond;
     layer1_node12_MUX_bit_math_h_l860_c3_f017_iftrue <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_iftrue;
     layer1_node12_MUX_bit_math_h_l860_c3_f017_iffalse <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_iffalse;
     -- Outputs
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_return_output := layer1_node12_MUX_bit_math_h_l860_c3_f017_return_output;

     -- layer1_node27_MUX[bit_math_h_l1025_c3_7ac4] LATENCY=0
     -- Inputs
     layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_cond <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_cond;
     layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iftrue <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iftrue;
     layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iffalse <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_iffalse;
     -- Outputs
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_return_output := layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_return_output;

     -- layer1_node18_MUX[bit_math_h_l926_c3_ab1a] LATENCY=0
     -- Inputs
     layer1_node18_MUX_bit_math_h_l926_c3_ab1a_cond <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_cond;
     layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iftrue <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iftrue;
     layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iffalse <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_iffalse;
     -- Outputs
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_return_output := layer1_node18_MUX_bit_math_h_l926_c3_ab1a_return_output;

     -- layer1_node31_MUX[bit_math_h_l1069_c3_fc71] LATENCY=0
     -- Inputs
     layer1_node31_MUX_bit_math_h_l1069_c3_fc71_cond <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_cond;
     layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iftrue <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iftrue;
     layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iffalse <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_iffalse;
     -- Outputs
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_return_output := layer1_node31_MUX_bit_math_h_l1069_c3_fc71_return_output;

     -- layer1_node8_MUX[bit_math_h_l816_c3_7279] LATENCY=0
     -- Inputs
     layer1_node8_MUX_bit_math_h_l816_c3_7279_cond <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_cond;
     layer1_node8_MUX_bit_math_h_l816_c3_7279_iftrue <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_iftrue;
     layer1_node8_MUX_bit_math_h_l816_c3_7279_iffalse <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_iffalse;
     -- Outputs
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_return_output := layer1_node8_MUX_bit_math_h_l816_c3_7279_return_output;

     -- layer1_node10_MUX[bit_math_h_l838_c3_e624] LATENCY=0
     -- Inputs
     layer1_node10_MUX_bit_math_h_l838_c3_e624_cond <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_cond;
     layer1_node10_MUX_bit_math_h_l838_c3_e624_iftrue <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_iftrue;
     layer1_node10_MUX_bit_math_h_l838_c3_e624_iffalse <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_iffalse;
     -- Outputs
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_return_output := layer1_node10_MUX_bit_math_h_l838_c3_e624_return_output;

     -- layer1_node6_MUX[bit_math_h_l794_c3_59a7] LATENCY=0
     -- Inputs
     layer1_node6_MUX_bit_math_h_l794_c3_59a7_cond <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_cond;
     layer1_node6_MUX_bit_math_h_l794_c3_59a7_iftrue <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_iftrue;
     layer1_node6_MUX_bit_math_h_l794_c3_59a7_iffalse <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_iffalse;
     -- Outputs
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_return_output := layer1_node6_MUX_bit_math_h_l794_c3_59a7_return_output;

     -- layer1_node0_MUX[bit_math_h_l728_c3_67cd] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l728_c3_67cd_cond <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_cond;
     layer1_node0_MUX_bit_math_h_l728_c3_67cd_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_iftrue;
     layer1_node0_MUX_bit_math_h_l728_c3_67cd_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_return_output := layer1_node0_MUX_bit_math_h_l728_c3_67cd_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iffalse := VAR_layer1_node0_MUX_bit_math_h_l728_c3_67cd_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iffalse := VAR_layer1_node10_MUX_bit_math_h_l838_c3_e624_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iftrue := VAR_layer1_node11_MUX_bit_math_h_l849_c3_0669_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_iffalse := VAR_layer1_node12_MUX_bit_math_h_l860_c3_f017_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_iftrue := VAR_layer1_node13_MUX_bit_math_h_l871_c3_9f0e_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iffalse := VAR_layer1_node14_MUX_bit_math_h_l882_c3_9be0_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iftrue := VAR_layer1_node15_MUX_bit_math_h_l893_c3_db88_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_iffalse := VAR_layer1_node16_MUX_bit_math_h_l904_c3_fdb3_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_iftrue := VAR_layer1_node17_MUX_bit_math_h_l915_c3_bba5_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iffalse := VAR_layer1_node18_MUX_bit_math_h_l926_c3_ab1a_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iftrue := VAR_layer1_node19_MUX_bit_math_h_l937_c3_1a24_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iftrue := VAR_layer1_node1_MUX_bit_math_h_l739_c3_5e54_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iffalse := VAR_layer1_node20_MUX_bit_math_h_l948_c3_2dbc_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iftrue := VAR_layer1_node21_MUX_bit_math_h_l959_c3_f718_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_iffalse := VAR_layer1_node22_MUX_bit_math_h_l970_c3_3aa5_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_iftrue := VAR_layer1_node23_MUX_bit_math_h_l981_c3_d2b9_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iffalse := VAR_layer1_node24_MUX_bit_math_h_l992_c3_8792_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iftrue := VAR_layer1_node25_MUX_bit_math_h_l1003_c3_2c90_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iffalse := VAR_layer1_node26_MUX_bit_math_h_l1014_c3_f8c1_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iftrue := VAR_layer1_node27_MUX_bit_math_h_l1025_c3_7ac4_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iffalse := VAR_layer1_node28_MUX_bit_math_h_l1036_c3_deef_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iftrue := VAR_layer1_node29_MUX_bit_math_h_l1047_c3_d4d6_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iffalse := VAR_layer1_node2_MUX_bit_math_h_l750_c3_386d_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iffalse := VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d1f5_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iftrue := VAR_layer1_node31_MUX_bit_math_h_l1069_c3_fc71_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iftrue := VAR_layer1_node3_MUX_bit_math_h_l761_c3_c96d_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_iffalse := VAR_layer1_node4_MUX_bit_math_h_l772_c3_535b_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_iftrue := VAR_layer1_node5_MUX_bit_math_h_l783_c3_7132_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iffalse := VAR_layer1_node6_MUX_bit_math_h_l794_c3_59a7_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iftrue := VAR_layer1_node7_MUX_bit_math_h_l805_c3_a7b7_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iffalse := VAR_layer1_node8_MUX_bit_math_h_l816_c3_7279_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iftrue := VAR_layer1_node9_MUX_bit_math_h_l827_c3_90fc_return_output;
     -- layer2_node7_MUX[bit_math_h_l1163_c3_d44d] LATENCY=0
     -- Inputs
     layer2_node7_MUX_bit_math_h_l1163_c3_d44d_cond <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_cond;
     layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iftrue <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iftrue;
     layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iffalse <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_iffalse;
     -- Outputs
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_return_output := layer2_node7_MUX_bit_math_h_l1163_c3_d44d_return_output;

     -- layer2_node13_MUX[bit_math_h_l1229_c3_d88d] LATENCY=0
     -- Inputs
     layer2_node13_MUX_bit_math_h_l1229_c3_d88d_cond <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_cond;
     layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iftrue <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iftrue;
     layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iffalse <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_iffalse;
     -- Outputs
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_return_output := layer2_node13_MUX_bit_math_h_l1229_c3_d88d_return_output;

     -- layer2_node3_MUX[bit_math_h_l1119_c3_b25e] LATENCY=0
     -- Inputs
     layer2_node3_MUX_bit_math_h_l1119_c3_b25e_cond <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_cond;
     layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iftrue <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iftrue;
     layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iffalse <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_iffalse;
     -- Outputs
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_return_output := layer2_node3_MUX_bit_math_h_l1119_c3_b25e_return_output;

     -- layer2_node2_MUX[bit_math_h_l1108_c3_922a] LATENCY=0
     -- Inputs
     layer2_node2_MUX_bit_math_h_l1108_c3_922a_cond <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_cond;
     layer2_node2_MUX_bit_math_h_l1108_c3_922a_iftrue <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_iftrue;
     layer2_node2_MUX_bit_math_h_l1108_c3_922a_iffalse <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_iffalse;
     -- Outputs
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_return_output := layer2_node2_MUX_bit_math_h_l1108_c3_922a_return_output;

     -- layer2_node6_MUX[bit_math_h_l1152_c3_d917] LATENCY=0
     -- Inputs
     layer2_node6_MUX_bit_math_h_l1152_c3_d917_cond <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_cond;
     layer2_node6_MUX_bit_math_h_l1152_c3_d917_iftrue <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_iftrue;
     layer2_node6_MUX_bit_math_h_l1152_c3_d917_iffalse <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_iffalse;
     -- Outputs
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_return_output := layer2_node6_MUX_bit_math_h_l1152_c3_d917_return_output;

     -- layer2_node4_MUX[bit_math_h_l1130_c3_5fd5] LATENCY=0
     -- Inputs
     layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_cond <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_cond;
     layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iftrue <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iftrue;
     layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iffalse <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_iffalse;
     -- Outputs
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_return_output := layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_return_output;

     -- layer2_node10_MUX[bit_math_h_l1196_c3_c6ad] LATENCY=0
     -- Inputs
     layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_cond <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_cond;
     layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iftrue <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iftrue;
     layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iffalse <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_iffalse;
     -- Outputs
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_return_output := layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_return_output;

     -- layer2_node0_MUX[bit_math_h_l1086_c3_5a52] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l1086_c3_5a52_cond <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_cond;
     layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iftrue;
     layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_return_output := layer2_node0_MUX_bit_math_h_l1086_c3_5a52_return_output;

     -- layer2_node1_MUX[bit_math_h_l1097_c3_fc1c] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_cond <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_cond;
     layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iftrue;
     layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_return_output := layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_return_output;

     -- layer2_node5_MUX[bit_math_h_l1141_c3_6ecd] LATENCY=0
     -- Inputs
     layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_cond <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_cond;
     layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iftrue <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iftrue;
     layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iffalse <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_iffalse;
     -- Outputs
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_return_output := layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_return_output;

     -- layer2_node11_MUX[bit_math_h_l1207_c3_e593] LATENCY=0
     -- Inputs
     layer2_node11_MUX_bit_math_h_l1207_c3_e593_cond <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_cond;
     layer2_node11_MUX_bit_math_h_l1207_c3_e593_iftrue <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_iftrue;
     layer2_node11_MUX_bit_math_h_l1207_c3_e593_iffalse <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_iffalse;
     -- Outputs
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_return_output := layer2_node11_MUX_bit_math_h_l1207_c3_e593_return_output;

     -- layer2_node14_MUX[bit_math_h_l1240_c3_d3d6] LATENCY=0
     -- Inputs
     layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_cond <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_cond;
     layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iftrue <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iftrue;
     layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iffalse <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_iffalse;
     -- Outputs
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_return_output := layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_return_output;

     -- layer2_node8_MUX[bit_math_h_l1174_c3_d504] LATENCY=0
     -- Inputs
     layer2_node8_MUX_bit_math_h_l1174_c3_d504_cond <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_cond;
     layer2_node8_MUX_bit_math_h_l1174_c3_d504_iftrue <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_iftrue;
     layer2_node8_MUX_bit_math_h_l1174_c3_d504_iffalse <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_iffalse;
     -- Outputs
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_return_output := layer2_node8_MUX_bit_math_h_l1174_c3_d504_return_output;

     -- layer2_node15_MUX[bit_math_h_l1251_c3_03ac] LATENCY=0
     -- Inputs
     layer2_node15_MUX_bit_math_h_l1251_c3_03ac_cond <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_cond;
     layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iftrue <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iftrue;
     layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iffalse <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_iffalse;
     -- Outputs
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_return_output := layer2_node15_MUX_bit_math_h_l1251_c3_03ac_return_output;

     -- layer2_node12_MUX[bit_math_h_l1218_c3_ed0c] LATENCY=0
     -- Inputs
     layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_cond <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_cond;
     layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iftrue <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iftrue;
     layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iffalse <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_iffalse;
     -- Outputs
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_return_output := layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_return_output;

     -- layer2_node9_MUX[bit_math_h_l1185_c3_8a90] LATENCY=0
     -- Inputs
     layer2_node9_MUX_bit_math_h_l1185_c3_8a90_cond <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_cond;
     layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iftrue <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iftrue;
     layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iffalse <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_iffalse;
     -- Outputs
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_return_output := layer2_node9_MUX_bit_math_h_l1185_c3_8a90_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_iffalse := VAR_layer2_node0_MUX_bit_math_h_l1086_c3_5a52_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iffalse := VAR_layer2_node10_MUX_bit_math_h_l1196_c3_c6ad_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iftrue := VAR_layer2_node11_MUX_bit_math_h_l1207_c3_e593_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iffalse := VAR_layer2_node12_MUX_bit_math_h_l1218_c3_ed0c_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iftrue := VAR_layer2_node13_MUX_bit_math_h_l1229_c3_d88d_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_iffalse := VAR_layer2_node14_MUX_bit_math_h_l1240_c3_d3d6_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_iftrue := VAR_layer2_node15_MUX_bit_math_h_l1251_c3_03ac_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_iftrue := VAR_layer2_node1_MUX_bit_math_h_l1097_c3_fc1c_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_iffalse := VAR_layer2_node2_MUX_bit_math_h_l1108_c3_922a_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_iftrue := VAR_layer2_node3_MUX_bit_math_h_l1119_c3_b25e_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_iffalse := VAR_layer2_node4_MUX_bit_math_h_l1130_c3_5fd5_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_iftrue := VAR_layer2_node5_MUX_bit_math_h_l1141_c3_6ecd_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iffalse := VAR_layer2_node6_MUX_bit_math_h_l1152_c3_d917_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iftrue := VAR_layer2_node7_MUX_bit_math_h_l1163_c3_d44d_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_iffalse := VAR_layer2_node8_MUX_bit_math_h_l1174_c3_d504_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_iftrue := VAR_layer2_node9_MUX_bit_math_h_l1185_c3_8a90_return_output;
     -- layer3_node0_MUX[bit_math_h_l1268_c3_6917] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l1268_c3_6917_cond <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_cond;
     layer3_node0_MUX_bit_math_h_l1268_c3_6917_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_iftrue;
     layer3_node0_MUX_bit_math_h_l1268_c3_6917_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_return_output := layer3_node0_MUX_bit_math_h_l1268_c3_6917_return_output;

     -- layer3_node3_MUX[bit_math_h_l1301_c3_fb21] LATENCY=0
     -- Inputs
     layer3_node3_MUX_bit_math_h_l1301_c3_fb21_cond <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_cond;
     layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iftrue <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iftrue;
     layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iffalse <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_iffalse;
     -- Outputs
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_return_output := layer3_node3_MUX_bit_math_h_l1301_c3_fb21_return_output;

     -- layer3_node4_MUX[bit_math_h_l1312_c3_f274] LATENCY=0
     -- Inputs
     layer3_node4_MUX_bit_math_h_l1312_c3_f274_cond <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_cond;
     layer3_node4_MUX_bit_math_h_l1312_c3_f274_iftrue <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_iftrue;
     layer3_node4_MUX_bit_math_h_l1312_c3_f274_iffalse <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_iffalse;
     -- Outputs
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_return_output := layer3_node4_MUX_bit_math_h_l1312_c3_f274_return_output;

     -- layer3_node7_MUX[bit_math_h_l1345_c3_969c] LATENCY=0
     -- Inputs
     layer3_node7_MUX_bit_math_h_l1345_c3_969c_cond <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_cond;
     layer3_node7_MUX_bit_math_h_l1345_c3_969c_iftrue <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_iftrue;
     layer3_node7_MUX_bit_math_h_l1345_c3_969c_iffalse <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_iffalse;
     -- Outputs
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_return_output := layer3_node7_MUX_bit_math_h_l1345_c3_969c_return_output;

     -- layer3_node6_MUX[bit_math_h_l1334_c3_41a0] LATENCY=0
     -- Inputs
     layer3_node6_MUX_bit_math_h_l1334_c3_41a0_cond <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_cond;
     layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iftrue <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iftrue;
     layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iffalse <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_iffalse;
     -- Outputs
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_return_output := layer3_node6_MUX_bit_math_h_l1334_c3_41a0_return_output;

     -- layer3_node5_MUX[bit_math_h_l1323_c3_6b46] LATENCY=0
     -- Inputs
     layer3_node5_MUX_bit_math_h_l1323_c3_6b46_cond <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_cond;
     layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iftrue <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iftrue;
     layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iffalse <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_iffalse;
     -- Outputs
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_return_output := layer3_node5_MUX_bit_math_h_l1323_c3_6b46_return_output;

     -- layer3_node2_MUX[bit_math_h_l1290_c3_769c] LATENCY=0
     -- Inputs
     layer3_node2_MUX_bit_math_h_l1290_c3_769c_cond <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_cond;
     layer3_node2_MUX_bit_math_h_l1290_c3_769c_iftrue <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_iftrue;
     layer3_node2_MUX_bit_math_h_l1290_c3_769c_iffalse <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_iffalse;
     -- Outputs
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_return_output := layer3_node2_MUX_bit_math_h_l1290_c3_769c_return_output;

     -- layer3_node1_MUX[bit_math_h_l1279_c3_e270] LATENCY=0
     -- Inputs
     layer3_node1_MUX_bit_math_h_l1279_c3_e270_cond <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_cond;
     layer3_node1_MUX_bit_math_h_l1279_c3_e270_iftrue <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_iftrue;
     layer3_node1_MUX_bit_math_h_l1279_c3_e270_iffalse <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_iffalse;
     -- Outputs
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_return_output := layer3_node1_MUX_bit_math_h_l1279_c3_e270_return_output;

     -- Submodule level 5
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iffalse := VAR_layer3_node0_MUX_bit_math_h_l1268_c3_6917_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iftrue := VAR_layer3_node1_MUX_bit_math_h_l1279_c3_e270_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iffalse := VAR_layer3_node2_MUX_bit_math_h_l1290_c3_769c_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iftrue := VAR_layer3_node3_MUX_bit_math_h_l1301_c3_fb21_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_iffalse := VAR_layer3_node4_MUX_bit_math_h_l1312_c3_f274_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_iftrue := VAR_layer3_node5_MUX_bit_math_h_l1323_c3_6b46_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iffalse := VAR_layer3_node6_MUX_bit_math_h_l1334_c3_41a0_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iftrue := VAR_layer3_node7_MUX_bit_math_h_l1345_c3_969c_return_output;
     -- layer4_node0_MUX[bit_math_h_l1362_c3_b41d] LATENCY=0
     -- Inputs
     layer4_node0_MUX_bit_math_h_l1362_c3_b41d_cond <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_cond;
     layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iftrue <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iftrue;
     layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iffalse <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_iffalse;
     -- Outputs
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_return_output := layer4_node0_MUX_bit_math_h_l1362_c3_b41d_return_output;

     -- layer4_node2_MUX[bit_math_h_l1384_c3_3339] LATENCY=0
     -- Inputs
     layer4_node2_MUX_bit_math_h_l1384_c3_3339_cond <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_cond;
     layer4_node2_MUX_bit_math_h_l1384_c3_3339_iftrue <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_iftrue;
     layer4_node2_MUX_bit_math_h_l1384_c3_3339_iffalse <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_iffalse;
     -- Outputs
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_return_output := layer4_node2_MUX_bit_math_h_l1384_c3_3339_return_output;

     -- layer4_node1_MUX[bit_math_h_l1373_c3_f2a6] LATENCY=0
     -- Inputs
     layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_cond <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_cond;
     layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iftrue <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iftrue;
     layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iffalse <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_iffalse;
     -- Outputs
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_return_output := layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_return_output;

     -- layer4_node3_MUX[bit_math_h_l1395_c3_b75d] LATENCY=0
     -- Inputs
     layer4_node3_MUX_bit_math_h_l1395_c3_b75d_cond <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_cond;
     layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iftrue <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iftrue;
     layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iffalse <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_iffalse;
     -- Outputs
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_return_output := layer4_node3_MUX_bit_math_h_l1395_c3_b75d_return_output;

     -- Submodule level 6
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iffalse := VAR_layer4_node0_MUX_bit_math_h_l1362_c3_b41d_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iftrue := VAR_layer4_node1_MUX_bit_math_h_l1373_c3_f2a6_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iffalse := VAR_layer4_node2_MUX_bit_math_h_l1384_c3_3339_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iftrue := VAR_layer4_node3_MUX_bit_math_h_l1395_c3_b75d_return_output;
     -- layer5_node1_MUX[bit_math_h_l1423_c3_1d22] LATENCY=0
     -- Inputs
     layer5_node1_MUX_bit_math_h_l1423_c3_1d22_cond <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_cond;
     layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iftrue <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iftrue;
     layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iffalse <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_iffalse;
     -- Outputs
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_return_output := layer5_node1_MUX_bit_math_h_l1423_c3_1d22_return_output;

     -- layer5_node0_MUX[bit_math_h_l1412_c3_5f1f] LATENCY=0
     -- Inputs
     layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_cond <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_cond;
     layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iftrue <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iftrue;
     layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iffalse <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_iffalse;
     -- Outputs
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_return_output := layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_return_output;

     -- Submodule level 7
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_iffalse := VAR_layer5_node0_MUX_bit_math_h_l1412_c3_5f1f_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_iftrue := VAR_layer5_node1_MUX_bit_math_h_l1423_c3_1d22_return_output;
     -- layer6_node0_MUX[bit_math_h_l1440_c3_247e] LATENCY=0
     -- Inputs
     layer6_node0_MUX_bit_math_h_l1440_c3_247e_cond <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_cond;
     layer6_node0_MUX_bit_math_h_l1440_c3_247e_iftrue <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_iftrue;
     layer6_node0_MUX_bit_math_h_l1440_c3_247e_iffalse <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_iffalse;
     -- Outputs
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_return_output := layer6_node0_MUX_bit_math_h_l1440_c3_247e_return_output;

     -- Submodule level 8
     VAR_return_output := VAR_layer6_node0_MUX_bit_math_h_l1440_c3_247e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
