-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity and2_0CLK_9159c4aa is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end and2_0CLK_9159c4aa;
architecture arch of and2_0CLK_9159c4aa is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l884_c6_eaab]
signal BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal n16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l884_c2_5e0e]
signal t16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l892_c11_80a5]
signal BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l892_c7_14f3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l892_c7_14f3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l892_c7_14f3]
signal result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l892_c7_14f3]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l892_c7_14f3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l892_c7_14f3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l892_c7_14f3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l892_c7_14f3]
signal n16_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l892_c7_14f3]
signal t16_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l895_c11_e4bd]
signal BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal n16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l895_c7_a8dc]
signal t16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l898_c30_eb97]
signal sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l900_c11_bc18]
signal BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l900_c7_4be0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l900_c7_4be0]
signal result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l900_c7_4be0]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l900_c7_4be0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l900_c7_4be0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l900_c7_4be0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l900_c7_4be0]
signal n16_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(15 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l905_c22_b23d]
signal BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_left : unsigned(15 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_right : unsigned(15 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l907_c11_4495]
signal BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l907_c7_75b9]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l907_c7_75b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l907_c7_75b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab
BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_left,
BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_right,
BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e
result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e
result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e
result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e
result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e
result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- n16_MUX_uxn_opcodes_h_l884_c2_5e0e
n16_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
n16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- t16_MUX_uxn_opcodes_h_l884_c2_5e0e
t16_MUX_uxn_opcodes_h_l884_c2_5e0e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond,
t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue,
t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse,
t16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5
BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_left,
BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_right,
BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3
result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3
result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3
result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3
result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3
result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- n16_MUX_uxn_opcodes_h_l892_c7_14f3
n16_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
n16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
n16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
n16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- t16_MUX_uxn_opcodes_h_l892_c7_14f3
t16_MUX_uxn_opcodes_h_l892_c7_14f3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l892_c7_14f3_cond,
t16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue,
t16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse,
t16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd
BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_left,
BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_right,
BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc
result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc
result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc
result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc
result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc
result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- n16_MUX_uxn_opcodes_h_l895_c7_a8dc
n16_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
n16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- t16_MUX_uxn_opcodes_h_l895_c7_a8dc
t16_MUX_uxn_opcodes_h_l895_c7_a8dc : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond,
t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue,
t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse,
t16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output);

-- sp_relative_shift_uxn_opcodes_h_l898_c30_eb97
sp_relative_shift_uxn_opcodes_h_l898_c30_eb97 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_ins,
sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_x,
sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_y,
sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18
BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_left,
BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_right,
BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0
result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0
result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_cond,
result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0
result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0
result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_return_output);

-- n16_MUX_uxn_opcodes_h_l900_c7_4be0
n16_MUX_uxn_opcodes_h_l900_c7_4be0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l900_c7_4be0_cond,
n16_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue,
n16_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse,
n16_MUX_uxn_opcodes_h_l900_c7_4be0_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d
BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d : entity work.BIN_OP_AND_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_left,
BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_right,
BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495
BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_left,
BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_right,
BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9
result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9
result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 n16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 t16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 n16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 t16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 n16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 t16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output,
 sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_return_output,
 n16_MUX_uxn_opcodes_h_l900_c7_4be0_return_output,
 BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l889_c3_d371 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_558a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l904_c3_4627 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l900_l884_l892_DUPLICATE_6841_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l900_l884_l892_l895_DUPLICATE_7145_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l884_l892_l895_DUPLICATE_4d01_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l884_l907_l892_l895_DUPLICATE_2118_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_e871_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_1141_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l900_l895_DUPLICATE_4ac4_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l913_l880_DUPLICATE_626a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l904_c3_4627 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l904_c3_4627;
     VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l889_c3_d371 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l889_c3_d371;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_558a := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_558a;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_right := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_e871 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_e871_return_output := result.is_stack_operation_16bit;

     -- BIN_OP_EQ[uxn_opcodes_h_l907_c11_4495] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_left;
     BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output := BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l884_l907_l892_l895_DUPLICATE_2118 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l884_l907_l892_l895_DUPLICATE_2118_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l884_l892_l895_DUPLICATE_4d01 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l884_l892_l895_DUPLICATE_4d01_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l884_c6_eaab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_left;
     BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output := BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l905_c22_b23d] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_left;
     BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_return_output := BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l900_l884_l892_l895_DUPLICATE_7145 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l900_l884_l892_l895_DUPLICATE_7145_return_output := result.u16_value;

     -- sp_relative_shift[uxn_opcodes_h_l898_c30_eb97] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_ins;
     sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_x <= VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_x;
     sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_y <= VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_return_output := sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l900_l895_DUPLICATE_4ac4 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l900_l895_DUPLICATE_4ac4_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_1141 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_1141_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l895_c11_e4bd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_left;
     BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output := BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l892_c11_80a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l900_l884_l892_DUPLICATE_6841 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l900_l884_l892_DUPLICATE_6841_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l900_c11_bc18] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_left;
     BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output := BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output;

     -- Submodule level 1
     VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l905_c22_b23d_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l884_c6_eaab_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l892_c11_80a5_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l895_c11_e4bd_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l900_c11_bc18_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l907_c11_4495_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l884_l892_l895_DUPLICATE_4d01_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l884_l892_l895_DUPLICATE_4d01_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l884_l892_l895_DUPLICATE_4d01_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l900_l884_l892_l895_DUPLICATE_7145_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l900_l884_l892_l895_DUPLICATE_7145_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l900_l884_l892_l895_DUPLICATE_7145_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l900_l884_l892_l895_DUPLICATE_7145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_1141_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_1141_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_1141_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_1141_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l900_l884_l892_DUPLICATE_6841_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l900_l884_l892_DUPLICATE_6841_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l900_l884_l892_DUPLICATE_6841_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_e871_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_e871_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_e871_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l900_l907_l892_l895_DUPLICATE_e871_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l884_l907_l892_l895_DUPLICATE_2118_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l884_l907_l892_l895_DUPLICATE_2118_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l884_l907_l892_l895_DUPLICATE_2118_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l884_l907_l892_l895_DUPLICATE_2118_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l900_l895_DUPLICATE_4ac4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l900_l895_DUPLICATE_4ac4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l898_c30_eb97_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l900_c7_4be0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;

     -- t16_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := t16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l907_c7_75b9] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_return_output;

     -- n16_MUX[uxn_opcodes_h_l900_c7_4be0] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l900_c7_4be0_cond <= VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_cond;
     n16_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue;
     n16_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_return_output := n16_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l907_c7_75b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l900_c7_4be0] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_cond;
     result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_return_output := result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l907_c7_75b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l900_c7_4be0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;

     -- Submodule level 2
     VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := VAR_n16_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l907_c7_75b9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l907_c7_75b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l907_c7_75b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_t16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     -- n16_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := n16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l900_c7_4be0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;

     -- t16_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     t16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     t16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := t16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l900_c7_4be0] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l900_c7_4be0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_n16_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l900_c7_4be0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_t16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l895_c7_a8dc] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;

     -- t16_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := t16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- n16_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     n16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     n16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := n16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_n16_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l895_c7_a8dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- n16_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := n16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l892_c7_14f3] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l892_c7_14f3_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l884_c2_5e0e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l913_l880_DUPLICATE_626a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l913_l880_DUPLICATE_626a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l884_c2_5e0e_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l913_l880_DUPLICATE_626a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l913_l880_DUPLICATE_626a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
