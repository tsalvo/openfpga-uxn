-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity neq_0CLK_57104a4d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_57104a4d;
architecture arch of neq_0CLK_57104a4d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1317_c6_3c39]
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1317_c2_68e5]
signal n8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1317_c2_68e5]
signal t8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1317_c2_68e5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1317_c2_68e5]
signal result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1317_c2_68e5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1317_c2_68e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1317_c2_68e5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1317_c2_68e5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1322_c11_bd59]
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1322_c7_28a5]
signal n8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1322_c7_28a5]
signal t8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1322_c7_28a5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1322_c7_28a5]
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1322_c7_28a5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1322_c7_28a5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1322_c7_28a5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1322_c7_28a5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1325_c11_a977]
signal BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1325_c7_ae11]
signal n8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1325_c7_ae11]
signal t8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1325_c7_ae11]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1325_c7_ae11]
signal result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1325_c7_ae11]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1325_c7_ae11]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1325_c7_ae11]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1325_c7_ae11]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1329_c11_0ae9]
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1329_c7_a04d]
signal n8_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1329_c7_a04d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1329_c7_a04d]
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1329_c7_a04d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1329_c7_a04d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1329_c7_a04d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1329_c7_a04d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1332_c11_b195]
signal BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1332_c7_f093]
signal n8_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1332_c7_f093]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1332_c7_f093]
signal result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1332_c7_f093]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1332_c7_f093]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1332_c7_f093]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1332_c7_f093]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1335_c30_405b]
signal sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1338_c21_0ed6]
signal BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1338_c21_beb9]
signal MUX_uxn_opcodes_h_l1338_c21_beb9_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1338_c21_beb9_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1338_c21_beb9_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1338_c21_beb9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1340_c11_7d67]
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1340_c7_b6ba]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1340_c7_b6ba]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1340_c7_b6ba]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39
BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_left,
BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_right,
BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output);

-- n8_MUX_uxn_opcodes_h_l1317_c2_68e5
n8_MUX_uxn_opcodes_h_l1317_c2_68e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond,
n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue,
n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse,
n8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

-- t8_MUX_uxn_opcodes_h_l1317_c2_68e5
t8_MUX_uxn_opcodes_h_l1317_c2_68e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond,
t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue,
t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse,
t8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5
result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5
result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_left,
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_right,
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output);

-- n8_MUX_uxn_opcodes_h_l1322_c7_28a5
n8_MUX_uxn_opcodes_h_l1322_c7_28a5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond,
n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue,
n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse,
n8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output);

-- t8_MUX_uxn_opcodes_h_l1322_c7_28a5
t8_MUX_uxn_opcodes_h_l1322_c7_28a5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond,
t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue,
t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse,
t8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977
BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_left,
BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_right,
BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output);

-- n8_MUX_uxn_opcodes_h_l1325_c7_ae11
n8_MUX_uxn_opcodes_h_l1325_c7_ae11 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond,
n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue,
n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse,
n8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output);

-- t8_MUX_uxn_opcodes_h_l1325_c7_ae11
t8_MUX_uxn_opcodes_h_l1325_c7_ae11 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond,
t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue,
t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse,
t8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11
result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_cond,
result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11
result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11
result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11
result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11
result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_left,
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_right,
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output);

-- n8_MUX_uxn_opcodes_h_l1329_c7_a04d
n8_MUX_uxn_opcodes_h_l1329_c7_a04d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1329_c7_a04d_cond,
n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue,
n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse,
n8_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195
BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_left,
BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_right,
BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output);

-- n8_MUX_uxn_opcodes_h_l1332_c7_f093
n8_MUX_uxn_opcodes_h_l1332_c7_f093 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1332_c7_f093_cond,
n8_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue,
n8_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse,
n8_MUX_uxn_opcodes_h_l1332_c7_f093_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093
result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_cond,
result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1335_c30_405b
sp_relative_shift_uxn_opcodes_h_l1335_c30_405b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_ins,
sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_x,
sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_y,
sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6
BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_left,
BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_right,
BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_return_output);

-- MUX_uxn_opcodes_h_l1338_c21_beb9
MUX_uxn_opcodes_h_l1338_c21_beb9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1338_c21_beb9_cond,
MUX_uxn_opcodes_h_l1338_c21_beb9_iftrue,
MUX_uxn_opcodes_h_l1338_c21_beb9_iffalse,
MUX_uxn_opcodes_h_l1338_c21_beb9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67
BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_left,
BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_right,
BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output,
 n8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
 t8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output,
 n8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output,
 t8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output,
 n8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output,
 t8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output,
 n8_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output,
 n8_MUX_uxn_opcodes_h_l1332_c7_f093_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output,
 sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_return_output,
 MUX_uxn_opcodes_h_l1338_c21_beb9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1319_c3_3613 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1323_c3_602e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_b5db : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1330_c3_ec05 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1337_c3_25be : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1332_c7_f093_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_c6fd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_51ab_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_496e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_1b88_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1340_l1332_l1329_l1325_l1322_DUPLICATE_98dc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1346_l1313_DUPLICATE_eaaf_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1319_c3_3613 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1319_c3_3613;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1330_c3_ec05 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1330_c3_ec05;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1337_c3_25be := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1337_c3_25be;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_b5db := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_b5db;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1323_c3_602e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1323_c3_602e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1340_l1332_l1329_l1325_l1322_DUPLICATE_98dc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1340_l1332_l1329_l1325_l1322_DUPLICATE_98dc_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_c6fd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_c6fd_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_1b88 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_1b88_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1340_c11_7d67] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_left;
     BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output := BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1322_c11_bd59] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_left;
     BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output := BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1338_c21_0ed6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1332_c7_f093] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1332_c7_f093_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1317_c6_3c39] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_left;
     BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output := BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_496e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_496e_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1332_c11_b195] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_left;
     BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output := BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1329_c11_0ae9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1335_c30_405b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_ins;
     sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_x;
     sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_return_output := sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_51ab LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_51ab_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1325_c11_a977] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_left;
     BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output := BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1317_c6_3c39_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_bd59_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1325_c11_a977_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_0ae9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1332_c11_b195_return_output;
     VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1338_c21_0ed6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c11_7d67_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_496e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_496e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_496e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_496e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_496e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1340_l1332_l1329_l1325_l1322_DUPLICATE_98dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1340_l1332_l1329_l1325_l1322_DUPLICATE_98dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1340_l1332_l1329_l1325_l1322_DUPLICATE_98dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1340_l1332_l1329_l1325_l1322_DUPLICATE_98dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1340_l1332_l1329_l1325_l1322_DUPLICATE_98dc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_1b88_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_1b88_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_1b88_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_1b88_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_1b88_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_51ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_51ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_51ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_51ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1317_l1340_l1329_l1325_l1322_DUPLICATE_51ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_c6fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_c6fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_c6fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_c6fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1317_l1332_l1329_l1325_l1322_DUPLICATE_c6fd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1332_c7_f093_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1335_c30_405b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1332_c7_f093] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1340_c7_b6ba] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output;

     -- MUX[uxn_opcodes_h_l1338_c21_beb9] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1338_c21_beb9_cond <= VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_cond;
     MUX_uxn_opcodes_h_l1338_c21_beb9_iftrue <= VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_iftrue;
     MUX_uxn_opcodes_h_l1338_c21_beb9_iffalse <= VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_return_output := MUX_uxn_opcodes_h_l1338_c21_beb9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1332_c7_f093] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;

     -- t8_MUX[uxn_opcodes_h_l1325_c7_ae11] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond <= VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond;
     t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue;
     t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output := t8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1340_c7_b6ba] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output;

     -- n8_MUX[uxn_opcodes_h_l1332_c7_f093] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1332_c7_f093_cond <= VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_cond;
     n8_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue;
     n8_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_return_output := n8_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1340_c7_b6ba] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue := VAR_MUX_uxn_opcodes_h_l1338_c21_beb9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1340_c7_b6ba_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1332_c7_f093] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1329_c7_a04d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;

     -- t8_MUX[uxn_opcodes_h_l1322_c7_28a5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond;
     t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue;
     t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output := t8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1329_c7_a04d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1329_c7_a04d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_cond;
     n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue;
     n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output := n8_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1329_c7_a04d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1332_c7_f093] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1332_c7_f093] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_return_output := result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1332_c7_f093] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1332_c7_f093_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;
     -- n8_MUX[uxn_opcodes_h_l1325_c7_ae11] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond <= VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_cond;
     n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue;
     n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output := n8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;

     -- t8_MUX[uxn_opcodes_h_l1317_c2_68e5] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond <= VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond;
     t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue;
     t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output := t8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1329_c7_a04d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1329_c7_a04d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1325_c7_ae11] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1329_c7_a04d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1325_c7_ae11] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1329_c7_a04d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_a04d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1325_c7_ae11] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output := result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1325_c7_ae11] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;

     -- n8_MUX[uxn_opcodes_h_l1322_c7_28a5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_cond;
     n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue;
     n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output := n8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1325_c7_ae11] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1322_c7_28a5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1322_c7_28a5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1325_c7_ae11] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1325_c7_ae11_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1317_c2_68e5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1322_c7_28a5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1322_c7_28a5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1322_c7_28a5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1317_c2_68e5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1322_c7_28a5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1317_c2_68e5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_cond;
     n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue;
     n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output := n8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_28a5_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1317_c2_68e5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1317_c2_68e5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1317_c2_68e5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1317_c2_68e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1346_l1313_DUPLICATE_eaaf LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1346_l1313_DUPLICATE_eaaf_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1317_c2_68e5_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1346_l1313_DUPLICATE_eaaf_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l1346_l1313_DUPLICATE_eaaf_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
