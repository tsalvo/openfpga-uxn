-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 36
entity nip2_0CLK_1a2ef46d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_1a2ef46d;
architecture arch of nip2_0CLK_1a2ef46d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2197_c6_55c6]
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c2_7cf0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2210_c11_b18e]
signal BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2210_c7_0803]
signal t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2210_c7_0803]
signal t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2210_c7_0803]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2210_c7_0803]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2210_c7_0803]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2210_c7_0803]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2210_c7_0803]
signal result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2213_c11_17be]
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2213_c7_ccb5]
signal t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2213_c7_ccb5]
signal t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c7_ccb5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c7_ccb5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c7_ccb5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c7_ccb5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2213_c7_ccb5]
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2215_c30_ba09]
signal sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2220_c11_5307]
signal BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2220_c7_2673]
signal t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2220_c7_2673]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2220_c7_2673]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2220_c7_2673]
signal result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2220_c7_2673]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e848( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6
BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_left,
BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_right,
BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0
t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0
t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e
BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_left,
BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_right,
BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2210_c7_0803
t16_low_MUX_uxn_opcodes_h_l2210_c7_0803 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_cond,
t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue,
t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse,
t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2210_c7_0803
t16_high_MUX_uxn_opcodes_h_l2210_c7_0803 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_cond,
t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue,
t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse,
t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803
result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803
result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803
result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803
result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_cond,
result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be
BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_left,
BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_right,
BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5
t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond,
t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue,
t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse,
t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5
t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond,
t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue,
t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse,
t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5
result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09
sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_ins,
sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_x,
sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_y,
sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307
BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_left,
BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_right,
BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2220_c7_2673
t16_low_MUX_uxn_opcodes_h_l2220_c7_2673 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_cond,
t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue,
t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse,
t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673
result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673
result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_cond,
result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673
result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output,
 t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output,
 t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_return_output,
 t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output,
 t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output,
 t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output,
 sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output,
 t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2202_c3_2f0b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2207_c3_83be : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2211_c3_c23d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2217_c3_1fac : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_ee7b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2220_c7_2673_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2222_c3_9fa8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2210_l2197_l2220_DUPLICATE_ac04_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2210_l2213_DUPLICATE_e010_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2210_l2220_DUPLICATE_1687_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2210_l2213_l2220_DUPLICATE_c0f2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2193_l2228_DUPLICATE_7744_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2211_c3_c23d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2211_c3_c23d;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_ee7b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_ee7b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2207_c3_83be := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2207_c3_83be;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2217_c3_1fac := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2217_c3_1fac;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2202_c3_2f0b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2202_c3_2f0b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_right := to_unsigned(2, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2222_c3_9fa8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2222_c3_9fa8;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse := t16_high;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse := t16_low;
     -- BIN_OP_EQ[uxn_opcodes_h_l2220_c11_5307] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_left;
     BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output := BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output := result.is_ram_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2213_c11_17be] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_left;
     BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output := BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2197_c6_55c6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2210_l2213_l2220_DUPLICATE_c0f2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2210_l2213_l2220_DUPLICATE_c0f2_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2210_l2197_l2220_DUPLICATE_ac04 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2210_l2197_l2220_DUPLICATE_ac04_return_output := result.u8_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2220_c7_2673] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2220_c7_2673_return_output := result.stack_address_sp_offset;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output := result.is_pc_updated;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2210_l2220_DUPLICATE_1687 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2210_l2220_DUPLICATE_1687_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2215_c30_ba09] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_ins;
     sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_x;
     sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_return_output := sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2210_c11_b18e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2210_l2213_DUPLICATE_e010 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2210_l2213_DUPLICATE_e010_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2197_c6_55c6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2210_c11_b18e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c11_17be_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2220_c11_5307_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2210_l2220_DUPLICATE_1687_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2210_l2220_DUPLICATE_1687_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2210_l2213_l2220_DUPLICATE_c0f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2210_l2213_l2220_DUPLICATE_c0f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2210_l2213_l2220_DUPLICATE_c0f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2210_l2213_DUPLICATE_e010_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2210_l2213_DUPLICATE_e010_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2210_l2197_l2220_DUPLICATE_ac04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2210_l2197_l2220_DUPLICATE_ac04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2210_l2197_l2220_DUPLICATE_ac04_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2197_c2_7cf0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2220_c7_2673_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2215_c30_ba09_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2220_c7_2673] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2220_c7_2673] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2220_c7_2673] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_return_output := result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2213_c7_ccb5] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond;
     t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output := t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2220_c7_2673] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c7_ccb5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2220_c7_2673] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_cond;
     t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_return_output := t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2220_c7_2673_return_output;
     -- t16_high_MUX[uxn_opcodes_h_l2210_c7_0803] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_cond;
     t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_return_output := t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c7_ccb5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c7_ccb5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2213_c7_ccb5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2210_c7_0803] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c7_ccb5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2213_c7_ccb5] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_cond;
     t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output := t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2213_c7_ccb5_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2210_c7_0803] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_return_output := result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2210_c7_0803] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2210_c7_0803] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2210_c7_0803] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2210_c7_0803] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_cond;
     t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_return_output := t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2210_c7_0803_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2197_c2_7cf0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;

     -- Submodule level 5
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2193_l2228_DUPLICATE_7744 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2193_l2228_DUPLICATE_7744_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e848(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2197_c2_7cf0_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2193_l2228_DUPLICATE_7744_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2193_l2228_DUPLICATE_7744_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
