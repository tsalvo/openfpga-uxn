-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity swp_0CLK_faaf4b1a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_faaf4b1a;
architecture arch of swp_0CLK_faaf4b1a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2415_c6_df47]
signal BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2415_c1_e5a5]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2415_c2_315d]
signal t8_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2415_c2_315d]
signal n8_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2415_c2_315d]
signal result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2415_c2_315d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2415_c2_315d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2415_c2_315d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2415_c2_315d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2415_c2_315d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l2416_c3_6176[uxn_opcodes_h_l2416_c3_6176]
signal printf_uxn_opcodes_h_l2416_c3_6176_uxn_opcodes_h_l2416_c3_6176_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2420_c11_43d8]
signal BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2420_c7_b6ae]
signal t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2420_c7_b6ae]
signal n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2420_c7_b6ae]
signal result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2420_c7_b6ae]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2420_c7_b6ae]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2420_c7_b6ae]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2420_c7_b6ae]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2420_c7_b6ae]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2423_c11_3f19]
signal BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2423_c7_8b31]
signal t8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2423_c7_8b31]
signal n8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2423_c7_8b31]
signal result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2423_c7_8b31]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2423_c7_8b31]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2423_c7_8b31]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2423_c7_8b31]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2423_c7_8b31]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2426_c11_a0f5]
signal BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2426_c7_fbd7]
signal n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2426_c7_fbd7]
signal result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2426_c7_fbd7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2426_c7_fbd7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2426_c7_fbd7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2426_c7_fbd7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2426_c7_fbd7]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2429_c30_ef68]
signal sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2434_c11_8dc3]
signal BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2434_c7_e3b7]
signal result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2434_c7_e3b7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2434_c7_e3b7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2434_c7_e3b7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2434_c7_e3b7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_2980]
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_db51]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_db51]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47
BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_left,
BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_right,
BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_return_output);

-- t8_MUX_uxn_opcodes_h_l2415_c2_315d
t8_MUX_uxn_opcodes_h_l2415_c2_315d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2415_c2_315d_cond,
t8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue,
t8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse,
t8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

-- n8_MUX_uxn_opcodes_h_l2415_c2_315d
n8_MUX_uxn_opcodes_h_l2415_c2_315d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2415_c2_315d_cond,
n8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue,
n8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse,
n8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d
result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d
result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d
result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d
result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

-- printf_uxn_opcodes_h_l2416_c3_6176_uxn_opcodes_h_l2416_c3_6176
printf_uxn_opcodes_h_l2416_c3_6176_uxn_opcodes_h_l2416_c3_6176 : entity work.printf_uxn_opcodes_h_l2416_c3_6176_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2416_c3_6176_uxn_opcodes_h_l2416_c3_6176_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8
BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_left,
BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_right,
BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output);

-- t8_MUX_uxn_opcodes_h_l2420_c7_b6ae
t8_MUX_uxn_opcodes_h_l2420_c7_b6ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond,
t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue,
t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse,
t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output);

-- n8_MUX_uxn_opcodes_h_l2420_c7_b6ae
n8_MUX_uxn_opcodes_h_l2420_c7_b6ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond,
n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue,
n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse,
n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae
result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond,
result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae
result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19
BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_left,
BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_right,
BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output);

-- t8_MUX_uxn_opcodes_h_l2423_c7_8b31
t8_MUX_uxn_opcodes_h_l2423_c7_8b31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond,
t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue,
t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse,
t8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output);

-- n8_MUX_uxn_opcodes_h_l2423_c7_8b31
n8_MUX_uxn_opcodes_h_l2423_c7_8b31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond,
n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue,
n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse,
n8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31
result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_cond,
result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31
result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31
result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31
result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31
result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5
BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_left,
BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_right,
BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output);

-- n8_MUX_uxn_opcodes_h_l2426_c7_fbd7
n8_MUX_uxn_opcodes_h_l2426_c7_fbd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond,
n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue,
n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse,
n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7
result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7
result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7
result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7
result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7
result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68
sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_ins,
sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_x,
sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_y,
sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3
BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_left,
BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_right,
BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7
result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond,
result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_left,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_right,
BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_return_output,
 t8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
 n8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output,
 t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output,
 n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output,
 t8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output,
 n8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output,
 n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output,
 sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2417_c3_e623 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2416_c3_6176_uxn_opcodes_h_l2416_c3_6176_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2421_c3_68d9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2431_c3_13cf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2436_c3_23b1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_081a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_df77_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2434_l2423_l2420_l2415_l2439_DUPLICATE_11c5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2415_l2426_l2420_l2423_DUPLICATE_9aa2_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2434_l2426_l2423_l2420_l2439_DUPLICATE_f9b5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2434_l2423_DUPLICATE_5c39_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2444_l2411_DUPLICATE_703f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2421_c3_68d9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2421_c3_68d9;
     VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2417_c3_e623 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2417_c3_e623;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2436_c3_23b1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2436_c3_23b1;
     VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2431_c3_13cf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2431_c3_13cf;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2426_c11_a0f5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2423_c11_3f19] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_left;
     BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output := BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_081a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_081a_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l2429_c30_ef68] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_ins;
     sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_x;
     sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_return_output := sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_df77 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_df77_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2420_c11_43d8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2434_l2423_l2420_l2415_l2439_DUPLICATE_11c5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2434_l2423_l2420_l2415_l2439_DUPLICATE_11c5_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2415_l2426_l2420_l2423_DUPLICATE_9aa2 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2415_l2426_l2420_l2423_DUPLICATE_9aa2_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2434_l2426_l2423_l2420_l2439_DUPLICATE_f9b5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2434_l2426_l2423_l2420_l2439_DUPLICATE_f9b5_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2439_c11_2980] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_left;
     BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_return_output := BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2434_l2423_DUPLICATE_5c39 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2434_l2423_DUPLICATE_5c39_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2415_c6_df47] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_left;
     BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output := BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2434_c11_8dc3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2415_c6_df47_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2420_c11_43d8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2423_c11_3f19_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2426_c11_a0f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2434_c11_8dc3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2439_c11_2980_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2415_l2426_l2420_l2423_DUPLICATE_9aa2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2415_l2426_l2420_l2423_DUPLICATE_9aa2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2415_l2426_l2420_l2423_DUPLICATE_9aa2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2415_l2426_l2420_l2423_DUPLICATE_9aa2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2434_l2426_l2423_l2420_l2439_DUPLICATE_f9b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2434_l2426_l2423_l2420_l2439_DUPLICATE_f9b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2434_l2426_l2423_l2420_l2439_DUPLICATE_f9b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2434_l2426_l2423_l2420_l2439_DUPLICATE_f9b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2434_l2426_l2423_l2420_l2439_DUPLICATE_f9b5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_df77_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_df77_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_df77_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_df77_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2434_l2423_l2420_l2415_l2439_DUPLICATE_11c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2434_l2423_l2420_l2415_l2439_DUPLICATE_11c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2434_l2423_l2420_l2415_l2439_DUPLICATE_11c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2434_l2423_l2420_l2415_l2439_DUPLICATE_11c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2434_l2423_l2420_l2415_l2439_DUPLICATE_11c5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2434_l2423_DUPLICATE_5c39_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2434_l2423_DUPLICATE_5c39_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_081a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_081a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_081a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2415_l2420_l2434_l2423_DUPLICATE_081a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2429_c30_ef68_return_output;
     -- n8_MUX[uxn_opcodes_h_l2426_c7_fbd7] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond <= VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond;
     n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue;
     n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output := n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2434_c7_e3b7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2439_c7_db51] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2415_c1_e5a5] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_return_output;

     -- t8_MUX[uxn_opcodes_h_l2423_c7_8b31] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond <= VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond;
     t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue;
     t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output := t8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2434_c7_e3b7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2434_c7_e3b7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2426_c7_fbd7] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2439_c7_db51] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2416_c3_6176_uxn_opcodes_h_l2416_c3_6176_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2415_c1_e5a5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2439_c7_db51_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2439_c7_db51_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2426_c7_fbd7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;

     -- n8_MUX[uxn_opcodes_h_l2423_c7_8b31] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond <= VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_cond;
     n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue;
     n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output := n8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2423_c7_8b31] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2426_c7_fbd7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;

     -- t8_MUX[uxn_opcodes_h_l2420_c7_b6ae] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond <= VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond;
     t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue;
     t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output := t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2434_c7_e3b7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2426_c7_fbd7] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output := result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;

     -- printf_uxn_opcodes_h_l2416_c3_6176[uxn_opcodes_h_l2416_c3_6176] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2416_c3_6176_uxn_opcodes_h_l2416_c3_6176_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2416_c3_6176_uxn_opcodes_h_l2416_c3_6176_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2434_c7_e3b7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2434_c7_e3b7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2420_c7_b6ae] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2426_c7_fbd7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;

     -- t8_MUX[uxn_opcodes_h_l2415_c2_315d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2415_c2_315d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_cond;
     t8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue;
     t8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output := t8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2426_c7_fbd7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2423_c7_8b31] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2423_c7_8b31] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2423_c7_8b31] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output := result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;

     -- n8_MUX[uxn_opcodes_h_l2420_c7_b6ae] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond <= VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond;
     n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue;
     n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output := n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2426_c7_fbd7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2420_c7_b6ae] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2423_c7_8b31] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2420_c7_b6ae] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output := result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2415_c2_315d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2420_c7_b6ae] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2423_c7_8b31] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;

     -- n8_MUX[uxn_opcodes_h_l2415_c2_315d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2415_c2_315d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_cond;
     n8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue;
     n8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output := n8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2423_c7_8b31_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2415_c2_315d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2415_c2_315d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2415_c2_315d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2420_c7_b6ae] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2420_c7_b6ae] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2420_c7_b6ae_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2415_c2_315d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2415_c2_315d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2444_l2411_DUPLICATE_703f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2444_l2411_DUPLICATE_703f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2415_c2_315d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2415_c2_315d_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2444_l2411_DUPLICATE_703f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l2444_l2411_DUPLICATE_703f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
