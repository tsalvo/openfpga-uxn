-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_f770903f is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_f770903f;
architecture arch of sft_0CLK_f770903f is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2177_c6_36f7]
signal BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2177_c2_5fc2]
signal tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2177_c2_5fc2]
signal n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2177_c2_5fc2]
signal result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2177_c2_5fc2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2177_c2_5fc2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2177_c2_5fc2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2177_c2_5fc2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2177_c2_5fc2]
signal t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2184_c11_1645]
signal BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2184_c7_f7da]
signal tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2184_c7_f7da]
signal n8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2184_c7_f7da]
signal result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2184_c7_f7da]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2184_c7_f7da]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2184_c7_f7da]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2184_c7_f7da]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2184_c7_f7da]
signal t8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_801e]
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2187_c7_4b2f]
signal tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2187_c7_4b2f]
signal n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_4b2f]
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_4b2f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_4b2f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_4b2f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_4b2f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l2187_c7_4b2f]
signal t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_1dab]
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2190_c7_386a]
signal tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2190_c7_386a]
signal n8_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_386a]
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_386a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_386a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_386a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_386a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2193_c30_3a91]
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2194_c18_1487]
signal BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2194_c11_65c0]
signal BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2194_c34_ea22]
signal CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2194_c11_af4f]
signal BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2199_c11_59f0]
signal BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2199_c7_026b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2199_c7_026b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2199_c7_026b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7
BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_left,
BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_right,
BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2
tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond,
tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue,
tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse,
tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

-- n8_MUX_uxn_opcodes_h_l2177_c2_5fc2
n8_MUX_uxn_opcodes_h_l2177_c2_5fc2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond,
n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue,
n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse,
n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2
result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2
result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2
result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

-- t8_MUX_uxn_opcodes_h_l2177_c2_5fc2
t8_MUX_uxn_opcodes_h_l2177_c2_5fc2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond,
t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue,
t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse,
t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645
BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_left,
BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_right,
BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da
tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond,
tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue,
tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse,
tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output);

-- n8_MUX_uxn_opcodes_h_l2184_c7_f7da
n8_MUX_uxn_opcodes_h_l2184_c7_f7da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond,
n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue,
n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse,
n8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da
result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_cond,
result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da
result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da
result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da
result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output);

-- t8_MUX_uxn_opcodes_h_l2184_c7_f7da
t8_MUX_uxn_opcodes_h_l2184_c7_f7da : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond,
t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue,
t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse,
t8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_left,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_right,
BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f
tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond,
tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue,
tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse,
tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output);

-- n8_MUX_uxn_opcodes_h_l2187_c7_4b2f
n8_MUX_uxn_opcodes_h_l2187_c7_4b2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond,
n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue,
n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse,
n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output);

-- t8_MUX_uxn_opcodes_h_l2187_c7_4b2f
t8_MUX_uxn_opcodes_h_l2187_c7_4b2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond,
t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue,
t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse,
t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_left,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_right,
BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2190_c7_386a
tmp8_MUX_uxn_opcodes_h_l2190_c7_386a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_cond,
tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue,
tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse,
tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output);

-- n8_MUX_uxn_opcodes_h_l2190_c7_386a
n8_MUX_uxn_opcodes_h_l2190_c7_386a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2190_c7_386a_cond,
n8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue,
n8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse,
n8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91
sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_ins,
sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_x,
sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_y,
sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487
BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_left,
BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_right,
BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0
BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0 : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_left,
BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_right,
BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22
CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22 : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_x,
CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f
BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_left,
BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_right,
BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0
BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_left,
BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_right,
BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b
result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b
result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output,
 tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
 n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
 t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output,
 tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output,
 n8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output,
 t8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output,
 tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output,
 n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output,
 t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output,
 tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output,
 n8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_return_output,
 sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_return_output,
 CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2181_c3_ce8a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_fc99 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2196_c3_29a0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_b43a : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2184_l2187_l2177_l2190_DUPLICATE_6a23_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_50c2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_c79a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2190_DUPLICATE_8bc1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_d066_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2205_l2173_DUPLICATE_5326_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_fc99 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_fc99;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2181_c3_ce8a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2181_c3_ce8a;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_b43a := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2200_c3_b43a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_right := to_unsigned(3, 2);
     VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_right := to_unsigned(15, 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2196_c3_29a0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2196_c3_29a0;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse := tmp8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_d066 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_d066_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2199_c11_59f0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2177_c6_36f7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_left;
     BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output := BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_50c2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_50c2_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2190_c11_1dab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_left;
     BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output := BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2193_c30_3a91] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_ins;
     sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_x;
     sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_return_output := sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_c79a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_c79a_return_output := result.sp_relative_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l2194_c18_1487] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_left;
     BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_return_output := BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2184_l2187_l2177_l2190_DUPLICATE_6a23 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2184_l2187_l2177_l2190_DUPLICATE_6a23_return_output := result.u8_value;

     -- CONST_SR_4[uxn_opcodes_h_l2194_c34_ea22] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_return_output := CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2187_c11_801e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2190_DUPLICATE_8bc1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2190_DUPLICATE_8bc1_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2184_c11_1645] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_left;
     BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output := BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2194_c18_1487_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2177_c6_36f7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2184_c11_1645_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2187_c11_801e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2190_c11_1dab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2199_c11_59f0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_c79a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_c79a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_c79a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_c79a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2190_DUPLICATE_8bc1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2190_DUPLICATE_8bc1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2190_DUPLICATE_8bc1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2190_DUPLICATE_8bc1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_50c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_50c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_50c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2184_l2199_l2187_l2177_DUPLICATE_50c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_d066_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2187_l2190_DUPLICATE_d066_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2184_l2187_l2177_l2190_DUPLICATE_6a23_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2184_l2187_l2177_l2190_DUPLICATE_6a23_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2184_l2187_l2177_l2190_DUPLICATE_6a23_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2184_l2187_l2177_l2190_DUPLICATE_6a23_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_right := VAR_CONST_SR_4_uxn_opcodes_h_l2194_c34_ea22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2193_c30_3a91_return_output;
     -- n8_MUX[uxn_opcodes_h_l2190_c7_386a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2190_c7_386a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_cond;
     n8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue;
     n8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output := n8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2190_c7_386a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2194_c11_65c0] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_left;
     BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_return_output := BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2187_c7_4b2f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond;
     t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue;
     t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output := t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2199_c7_026b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2199_c7_026b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2199_c7_026b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2194_c11_65c0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2199_c7_026b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2199_c7_026b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2199_c7_026b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2190_c7_386a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2194_c11_af4f] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_left;
     BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_return_output := BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2187_c7_4b2f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2190_c7_386a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2184_c7_f7da] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond <= VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond;
     t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue;
     t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output := t8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2190_c7_386a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2187_c7_4b2f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond;
     n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue;
     n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output := n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2194_c11_af4f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2187_c7_4b2f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2190_c7_386a] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_cond;
     tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output := tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2184_c7_f7da] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond <= VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond;
     n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue;
     n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output := n8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2187_c7_4b2f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2184_c7_f7da] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2187_c7_4b2f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2190_c7_386a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2177_c2_5fc2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond;
     t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue;
     t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output := t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2190_c7_386a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2184_c7_f7da] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2184_c7_f7da] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2184_c7_f7da] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2187_c7_4b2f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2177_c2_5fc2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond <= VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond;
     n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue;
     n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output := n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2177_c2_5fc2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2187_c7_4b2f] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_cond;
     tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output := tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2187_c7_4b2f_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2177_c2_5fc2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2177_c2_5fc2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2177_c2_5fc2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2184_c7_f7da] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_cond;
     tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output := tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2184_c7_f7da] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output := result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2184_c7_f7da_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2177_c2_5fc2] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond;
     tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output := tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2177_c2_5fc2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2205_l2173_DUPLICATE_5326 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2205_l2173_DUPLICATE_5326_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2177_c2_5fc2_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2205_l2173_DUPLICATE_5326_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l2205_l2173_DUPLICATE_5326_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
