-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity eor_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_64d180f1;
architecture arch of eor_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1099_c6_b1e9]
signal BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1099_c2_d350]
signal n8_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1099_c2_d350]
signal t8_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1099_c2_d350]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1112_c11_9788]
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1112_c7_a687]
signal n8_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1112_c7_a687]
signal t8_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1112_c7_a687]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1112_c7_a687]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1112_c7_a687]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1112_c7_a687]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1112_c7_a687]
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1115_c11_8d90]
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1115_c7_bc41]
signal n8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1115_c7_bc41]
signal t8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1115_c7_bc41]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1115_c7_bc41]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1115_c7_bc41]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1115_c7_bc41]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1115_c7_bc41]
signal result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1118_c11_120c]
signal BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1118_c7_96ab]
signal n8_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1118_c7_96ab]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1118_c7_96ab]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1118_c7_96ab]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1118_c7_96ab]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1118_c7_96ab]
signal result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1120_c30_c71e]
signal sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1123_c21_6442]
signal BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e848( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9
BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_left,
BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_right,
BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output);

-- n8_MUX_uxn_opcodes_h_l1099_c2_d350
n8_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
n8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
n8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
n8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- t8_MUX_uxn_opcodes_h_l1099_c2_d350
t8_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
t8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
t8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
t8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_left,
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_right,
BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output);

-- n8_MUX_uxn_opcodes_h_l1112_c7_a687
n8_MUX_uxn_opcodes_h_l1112_c7_a687 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1112_c7_a687_cond,
n8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue,
n8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse,
n8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output);

-- t8_MUX_uxn_opcodes_h_l1112_c7_a687
t8_MUX_uxn_opcodes_h_l1112_c7_a687 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1112_c7_a687_cond,
t8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue,
t8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse,
t8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_cond,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90
BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_left,
BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_right,
BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output);

-- n8_MUX_uxn_opcodes_h_l1115_c7_bc41
n8_MUX_uxn_opcodes_h_l1115_c7_bc41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond,
n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue,
n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse,
n8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output);

-- t8_MUX_uxn_opcodes_h_l1115_c7_bc41
t8_MUX_uxn_opcodes_h_l1115_c7_bc41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond,
t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue,
t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse,
t8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_cond,
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c
BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_left,
BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_right,
BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output);

-- n8_MUX_uxn_opcodes_h_l1118_c7_96ab
n8_MUX_uxn_opcodes_h_l1118_c7_96ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1118_c7_96ab_cond,
n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue,
n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse,
n8_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_cond,
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e
sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_ins,
sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_x,
sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_y,
sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442
BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442 : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_left,
BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_right,
BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output,
 n8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 t8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output,
 n8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output,
 t8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output,
 n8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output,
 t8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output,
 n8_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output,
 sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1104_c3_df64 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1109_c3_1143 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1113_c3_0138 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1122_c3_8e56 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_578d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_8305_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_c7b9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_2ad1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_cc47_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1127_l1095_DUPLICATE_c740_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1104_c3_df64 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1104_c3_df64;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1109_c3_1143 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1109_c3_1143;
     VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1113_c3_0138 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1113_c3_0138;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1122_c3_8e56 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1122_c3_8e56;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1099_c6_b1e9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1120_c30_c71e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_ins;
     sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_x;
     sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_return_output := sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1112_c11_9788] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_left;
     BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output := BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_c7b9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_c7b9_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_578d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_578d_return_output := result.u8_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1099_c2_d350_return_output := result.is_stack_index_flipped;

     -- BIN_OP_XOR[uxn_opcodes_h_l1123_c21_6442] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_left;
     BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_return_output := BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_8305 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_8305_return_output := result.is_stack_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1099_c2_d350_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_cc47 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_cc47_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1118_c11_120c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_2ad1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_2ad1_return_output := result.is_opc_done;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1099_c2_d350_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1115_c11_8d90] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_left;
     BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output := BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1099_c2_d350_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1099_c6_b1e9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1112_c11_9788_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1115_c11_8d90_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1118_c11_120c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1123_c21_6442_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_c7b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_c7b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_c7b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_2ad1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_2ad1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_2ad1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_8305_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_8305_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1118_l1112_l1115_DUPLICATE_8305_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_cc47_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1118_l1115_DUPLICATE_cc47_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_578d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_578d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_578d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1099_l1118_l1112_l1115_DUPLICATE_578d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1099_c2_d350_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1099_c2_d350_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1099_c2_d350_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1099_c2_d350_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1120_c30_c71e_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- t8_MUX[uxn_opcodes_h_l1115_c7_bc41] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond <= VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond;
     t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue;
     t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output := t8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1118_c7_96ab] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;

     -- n8_MUX[uxn_opcodes_h_l1118_c7_96ab] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1118_c7_96ab_cond <= VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_cond;
     n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue;
     n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output := n8_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1118_c7_96ab] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1118_c7_96ab] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output := result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1118_c7_96ab] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1118_c7_96ab] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1118_c7_96ab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1115_c7_bc41] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1115_c7_bc41] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1115_c7_bc41] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output := result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;

     -- n8_MUX[uxn_opcodes_h_l1115_c7_bc41] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond <= VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_cond;
     n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue;
     n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output := n8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;

     -- t8_MUX[uxn_opcodes_h_l1112_c7_a687] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1112_c7_a687_cond <= VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_cond;
     t8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue;
     t8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output := t8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1115_c7_bc41] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1115_c7_bc41] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1115_c7_bc41_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;
     -- n8_MUX[uxn_opcodes_h_l1112_c7_a687] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1112_c7_a687_cond <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_cond;
     n8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue;
     n8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output := n8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1112_c7_a687] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1112_c7_a687] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;

     -- t8_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     t8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     t8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := t8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1112_c7_a687] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_return_output := result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1112_c7_a687] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1112_c7_a687] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1112_c7_a687_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- n8_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     n8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     n8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := n8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1099_c2_d350] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1099_c2_d350_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1127_l1095_DUPLICATE_c740 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1127_l1095_DUPLICATE_c740_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e848(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1099_c2_d350_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1099_c2_d350_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1127_l1095_DUPLICATE_c740_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l1127_l1095_DUPLICATE_c740_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
