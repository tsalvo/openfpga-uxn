-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity inc2_0CLK_180c5210 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_180c5210;
architecture arch of inc2_0CLK_180c5210 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1355_c6_9ffe]
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1355_c2_6bdb]
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1368_c11_f85d]
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1368_c7_9333]
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1368_c7_9333]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1368_c7_9333]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1368_c7_9333]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1368_c7_9333]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1368_c7_9333]
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1368_c7_9333]
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1371_c11_002d]
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1371_c7_de8c]
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1371_c7_de8c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1371_c7_de8c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1371_c7_de8c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1371_c7_de8c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1371_c7_de8c]
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1371_c7_de8c]
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1372_c13_bbde]
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_return_output : unsigned(8 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1373_c30_8184]
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_5303]
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c7_18b6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_18b6]
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_18b6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_18b6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1378_c7_18b6]
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1379_c37_54e2]
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1379_c37_4cbc]
signal MUX_uxn_opcodes_h_l1379_c37_4cbc_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_4cbc_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_4cbc_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1379_c37_4cbc_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1379_c14_7a9e]
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_922a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_opc_done := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_left,
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_right,
BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb
t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb
t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond,
t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue,
t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse,
t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_left,
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_right,
BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_cond,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1368_c7_9333
t16_high_MUX_uxn_opcodes_h_l1368_c7_9333 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_cond,
t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue,
t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse,
t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1368_c7_9333
t16_low_MUX_uxn_opcodes_h_l1368_c7_9333 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_cond,
t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue,
t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse,
t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_left,
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_right,
BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c
t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_cond,
t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue,
t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse,
t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c
t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_cond,
t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue,
t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse,
t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_left,
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_right,
BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1373_c30_8184
sp_relative_shift_uxn_opcodes_h_l1373_c30_8184 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_ins,
sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_x,
sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_y,
sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_left,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_right,
BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_cond,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6
t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_cond,
t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue,
t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse,
t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_left,
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_right,
BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_return_output);

-- MUX_uxn_opcodes_h_l1379_c37_4cbc
MUX_uxn_opcodes_h_l1379_c37_4cbc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1379_c37_4cbc_cond,
MUX_uxn_opcodes_h_l1379_c37_4cbc_iftrue,
MUX_uxn_opcodes_h_l1379_c37_4cbc_iffalse,
MUX_uxn_opcodes_h_l1379_c37_4cbc_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_left,
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_right,
BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_return_output,
 t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_return_output,
 t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output,
 t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output,
 t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_return_output,
 sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output,
 t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_return_output,
 MUX_uxn_opcodes_h_l1379_c37_4cbc_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_6d35 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_ed55 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_2c88 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_a012 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_uxn_opcodes_h_l1372_c3_5dde : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_return_output : unsigned(8 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_ef13 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_5e31 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_18b6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_uxn_opcodes_h_l1379_c3_762e : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_left : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c71_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_e6dd_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_d746_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_0c17_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1386_l1351_DUPLICATE_41cd_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_5e31 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1381_c3_5e31;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_2c88 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1369_c3_2c88;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_ed55 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1360_c3_ed55;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_6d35 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1365_c3_6d35;
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_ef13 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1380_c3_ef13;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_a012 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1375_c3_a012;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_left := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_left := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse := t16_high;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_left := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse := t16_low;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1378_c7_18b6] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_18b6_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1378_c11_5303] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_left;
     BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output := BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1379_c37_54e2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_d746 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_d746_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_0c17 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_0c17_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1371_c11_002d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1372_c13_bbde] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1355_c6_9ffe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_left;
     BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output := BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_e6dd LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_e6dd_return_output := result.sp_relative_shift;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c71 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c71_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l1373_c30_8184] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_ins;
     sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_x;
     sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_return_output := sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1368_c11_f85d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1355_c6_9ffe_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1368_c11_f85d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1371_c11_002d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c11_5303_return_output;
     VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1379_c37_54e2_return_output;
     VAR_t16_low_uxn_opcodes_h_l1372_c3_5dde := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1372_c13_bbde_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_e6dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1378_l1368_DUPLICATE_e6dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_d746_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_d746_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1371_l1378_l1368_DUPLICATE_d746_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_0c17_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1371_l1368_DUPLICATE_0c17_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c71_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c71_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1355_l1378_l1368_DUPLICATE_3c71_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1355_c2_6bdb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1378_c7_18b6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1373_c30_8184_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue := VAR_t16_low_uxn_opcodes_h_l1372_c3_5dde;
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue := VAR_t16_low_uxn_opcodes_h_l1372_c3_5dde;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1371_c7_de8c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- MUX[uxn_opcodes_h_l1379_c37_4cbc] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1379_c37_4cbc_cond <= VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_cond;
     MUX_uxn_opcodes_h_l1379_c37_4cbc_iftrue <= VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_iftrue;
     MUX_uxn_opcodes_h_l1379_c37_4cbc_iffalse <= VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_return_output := MUX_uxn_opcodes_h_l1379_c37_4cbc_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c7_18b6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1371_c7_de8c] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_cond;
     t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output := t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c7_18b6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c7_18b6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_right := VAR_MUX_uxn_opcodes_h_l1379_c37_4cbc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1371_c7_de8c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1371_c7_de8c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1368_c7_9333] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1368_c7_9333] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_cond;
     t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_return_output := t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1371_c7_de8c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1379_c14_7a9e] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_return_output;

     -- Submodule level 3
     VAR_t16_high_uxn_opcodes_h_l1379_c3_762e := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1379_c14_7a9e_return_output, 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue := VAR_t16_high_uxn_opcodes_h_l1379_c3_762e;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue := VAR_t16_high_uxn_opcodes_h_l1379_c3_762e;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1368_c7_9333] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1378_c7_18b6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output := result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1368_c7_9333] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1378_c7_18b6] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_cond;
     t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output := t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1368_c7_9333] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1378_c7_18b6_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1371_c7_de8c] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_cond;
     t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output := t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1371_c7_de8c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;

     -- Submodule level 5
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1371_c7_de8c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1368_c7_9333] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_return_output := result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1368_c7_9333] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_cond;
     t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_return_output := t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1368_c7_9333_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1355_c2_6bdb] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_cond;
     t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output := t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;

     -- Submodule level 7
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1386_l1351_DUPLICATE_41cd LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1386_l1351_DUPLICATE_41cd_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_922a(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1355_c2_6bdb_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1386_l1351_DUPLICATE_41cd_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l1386_l1351_DUPLICATE_41cd_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
