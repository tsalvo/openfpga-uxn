-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 46
entity jsr_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jsr_0CLK_fedec265;
architecture arch of jsr_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l754_c6_9e2c]
signal BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l754_c2_183f]
signal t8_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l754_c2_183f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l767_c11_af21]
signal BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l767_c7_b578]
signal t8_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l767_c7_b578]
signal result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l767_c7_b578]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l767_c7_b578]
signal result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l767_c7_b578]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l767_c7_b578]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l767_c7_b578]
signal result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l767_c7_b578]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l767_c7_b578]
signal result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l769_c30_d21a]
signal sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l771_c11_d4a7]
signal BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l771_c7_c39a]
signal t8_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l771_c7_c39a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l771_c7_c39a]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l771_c7_c39a]
signal result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l771_c7_c39a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l771_c7_c39a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l771_c7_c39a]
signal result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l771_c7_c39a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l771_c7_c39a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l779_c11_82b7]
signal BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l779_c7_a926]
signal result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l779_c7_a926]
signal result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l779_c7_a926]
signal result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l779_c7_a926]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l779_c7_a926]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l779_c7_a926]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(0 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l782_c31_e55a]
signal CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l784_c22_bb08]
signal BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_return_output : signed(17 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_1a75( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;
      base.is_pc_updated := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c
BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_left,
BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_right,
BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output);

-- t8_MUX_uxn_opcodes_h_l754_c2_183f
t8_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l754_c2_183f_cond,
t8_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
t8_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
t8_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f
result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f
result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21
BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_left,
BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_right,
BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output);

-- t8_MUX_uxn_opcodes_h_l767_c7_b578
t8_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l767_c7_b578_cond,
t8_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
t8_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
t8_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578
result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_cond,
result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578
result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_cond,
result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_return_output);

-- sp_relative_shift_uxn_opcodes_h_l769_c30_d21a
sp_relative_shift_uxn_opcodes_h_l769_c30_d21a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_ins,
sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_x,
sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_y,
sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7
BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_left,
BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_right,
BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output);

-- t8_MUX_uxn_opcodes_h_l771_c7_c39a
t8_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
t8_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
t8_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
t8_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a
result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a
result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7
BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_left,
BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_right,
BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926
result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_cond,
result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926
result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_cond,
result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_return_output);

-- CONST_SR_8_uxn_opcodes_h_l782_c31_e55a
CONST_SR_8_uxn_opcodes_h_l782_c31_e55a : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_x,
CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08
BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_left,
BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_right,
BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output,
 t8_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output,
 t8_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_return_output,
 sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output,
 t8_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_return_output,
 CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_9704 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_e5c9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l768_c3_d0b0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l774_c3_d097 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_7ec6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_73a4_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l784_c3_cb9e : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l780_c3_8263 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l779_c7_a926_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l781_c3_061b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l779_c7_a926_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l782_c21_0fa6_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l784_c27_e95e_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_return_output : signed(17 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l779_l767_l771_l754_DUPLICATE_7c93_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l779_l767_l754_DUPLICATE_33a5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_7df0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_10a3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_49f0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_dd3c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l788_l750_DUPLICATE_0aa4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_right := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l768_c3_d0b0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l768_c3_d0b0;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_9704 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l759_c3_9704;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l781_c3_061b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l781_c3_061b;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l774_c3_d097 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l774_c3_d097;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_e5c9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l764_c3_e5c9;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l780_c3_8263 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l780_c3_8263;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_7ec6 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l776_c3_7ec6;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_x := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_left := VAR_phase;
     VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_10a3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_10a3_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l771_c11_d4a7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_left;
     BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output := BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;

     -- CAST_TO_int8_t[uxn_opcodes_h_l784_c27_e95e] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l784_c27_e95e_return_output := CAST_TO_int8_t_uint8_t(
     t8);

     -- BIN_OP_EQ[uxn_opcodes_h_l779_c11_82b7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_left;
     BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output := BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l754_c6_9e2c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_left;
     BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output := BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l754_c2_183f_return_output := result.is_ram_write;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l777_c21_73a4] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_73a4_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_pc);

     -- CONST_SR_8[uxn_opcodes_h_l782_c31_e55a] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_x <= VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_return_output := CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l779_c7_a926] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l779_c7_a926_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_dd3c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_dd3c_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_7df0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_7df0_return_output := result.is_opc_done;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l779_c7_a926] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l779_c7_a926_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l779_l767_l754_DUPLICATE_33a5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l779_l767_l754_DUPLICATE_33a5_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l769_c30_d21a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_ins;
     sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_x;
     sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_return_output := sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l754_c2_183f_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l767_c11_af21] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_left;
     BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output := BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l779_l767_l771_l754_DUPLICATE_7c93 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l779_l767_l771_l754_DUPLICATE_7c93_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_49f0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_49f0_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l754_c6_9e2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l767_c11_af21_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l771_c11_d4a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l779_c11_82b7_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l784_c27_e95e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l777_c21_73a4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l779_l767_l771_l754_DUPLICATE_7c93_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l779_l767_l771_l754_DUPLICATE_7c93_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l779_l767_l771_l754_DUPLICATE_7c93_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l779_l767_l771_l754_DUPLICATE_7c93_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_7df0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_7df0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_7df0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_49f0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_49f0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l779_l767_l771_DUPLICATE_49f0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_10a3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_10a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_dd3c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l767_l771_DUPLICATE_dd3c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l779_l767_l754_DUPLICATE_33a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l779_l767_l754_DUPLICATE_33a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l779_l767_l754_DUPLICATE_33a5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l754_c2_183f_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l754_c2_183f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l779_c7_a926_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l779_c7_a926_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l769_c30_d21a_return_output;
     -- BIN_OP_PLUS[uxn_opcodes_h_l784_c22_bb08] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_left;
     BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_return_output := BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l782_c21_0fa6] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l782_c21_0fa6_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l782_c31_e55a_return_output);

     -- result_is_ram_write_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- t8_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     t8_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     t8_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := t8_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l779_c7_a926] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l779_c7_a926] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l779_c7_a926] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l779_c7_a926] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l784_c3_cb9e := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l784_c22_bb08_return_output)),16);
     VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l782_c21_0fa6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l779_c7_a926_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l779_c7_a926_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l779_c7_a926_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l779_c7_a926_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_t8_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue := VAR_result_u16_value_uxn_opcodes_h_l784_c3_cb9e;
     -- result_u16_value_MUX[uxn_opcodes_h_l779_c7_a926] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_cond;
     result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output := result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l779_c7_a926] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_cond;
     result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output := result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- t8_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     t8_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     t8_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_return_output := t8_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l779_c7_a926_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- t8_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     t8_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     t8_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_return_output := t8_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l771_c7_c39a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output := result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l771_c7_c39a_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l754_c2_183f_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output := result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l767_c7_b578] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_cond;
     result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output := result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l767_c7_b578_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l754_c2_183f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output := result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l788_l750_DUPLICATE_0aa4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l788_l750_DUPLICATE_0aa4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_1a75(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l754_c2_183f_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l754_c2_183f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l788_l750_DUPLICATE_0aa4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_1a75_uxn_opcodes_h_l788_l750_DUPLICATE_0aa4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
