-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity neq_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_6d7675a8;
architecture arch of neq_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1319_c6_a5f2]
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1319_c1_46a0]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1319_c2_d110]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1319_c2_d110]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1319_c2_d110]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1319_c2_d110]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1319_c2_d110]
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1319_c2_d110]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1319_c2_d110]
signal t8_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1319_c2_d110]
signal n8_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1320_c3_453d[uxn_opcodes_h_l1320_c3_453d]
signal printf_uxn_opcodes_h_l1320_c3_453d_uxn_opcodes_h_l1320_c3_453d_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1324_c11_2a30]
signal BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1324_c7_c247]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1324_c7_c247]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1324_c7_c247]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1324_c7_c247]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1324_c7_c247]
signal result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1324_c7_c247]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1324_c7_c247]
signal t8_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1324_c7_c247]
signal n8_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1327_c11_a578]
signal BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1327_c7_f738]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1327_c7_f738]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1327_c7_f738]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1327_c7_f738]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1327_c7_f738]
signal result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1327_c7_f738]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1327_c7_f738]
signal t8_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1327_c7_f738]
signal n8_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1331_c11_c290]
signal BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1331_c7_42b1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1331_c7_42b1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1331_c7_42b1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1331_c7_42b1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1331_c7_42b1]
signal result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1331_c7_42b1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1331_c7_42b1]
signal n8_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1334_c11_0023]
signal BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1334_c7_b2ef]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1334_c7_b2ef]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1334_c7_b2ef]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1334_c7_b2ef]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1334_c7_b2ef]
signal result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1334_c7_b2ef]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1334_c7_b2ef]
signal n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1337_c30_762f]
signal sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1340_c21_0dce]
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1340_c21_7540]
signal MUX_uxn_opcodes_h_l1340_c21_7540_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1340_c21_7540_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1340_c21_7540_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1340_c21_7540_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1342_c11_9c4c]
signal BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1342_c7_7f0c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1342_c7_7f0c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1342_c7_7f0c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2
BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_left,
BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_right,
BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110
result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_cond,
result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

-- t8_MUX_uxn_opcodes_h_l1319_c2_d110
t8_MUX_uxn_opcodes_h_l1319_c2_d110 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1319_c2_d110_cond,
t8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue,
t8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse,
t8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

-- n8_MUX_uxn_opcodes_h_l1319_c2_d110
n8_MUX_uxn_opcodes_h_l1319_c2_d110 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1319_c2_d110_cond,
n8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue,
n8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse,
n8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

-- printf_uxn_opcodes_h_l1320_c3_453d_uxn_opcodes_h_l1320_c3_453d
printf_uxn_opcodes_h_l1320_c3_453d_uxn_opcodes_h_l1320_c3_453d : entity work.printf_uxn_opcodes_h_l1320_c3_453d_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1320_c3_453d_uxn_opcodes_h_l1320_c3_453d_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30
BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_left,
BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_right,
BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247
result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247
result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247
result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247
result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_cond,
result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247
result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output);

-- t8_MUX_uxn_opcodes_h_l1324_c7_c247
t8_MUX_uxn_opcodes_h_l1324_c7_c247 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1324_c7_c247_cond,
t8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue,
t8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse,
t8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output);

-- n8_MUX_uxn_opcodes_h_l1324_c7_c247
n8_MUX_uxn_opcodes_h_l1324_c7_c247 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1324_c7_c247_cond,
n8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue,
n8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse,
n8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578
BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_left,
BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_right,
BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738
result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738
result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_cond,
result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output);

-- t8_MUX_uxn_opcodes_h_l1327_c7_f738
t8_MUX_uxn_opcodes_h_l1327_c7_f738 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1327_c7_f738_cond,
t8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue,
t8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse,
t8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output);

-- n8_MUX_uxn_opcodes_h_l1327_c7_f738
n8_MUX_uxn_opcodes_h_l1327_c7_f738 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1327_c7_f738_cond,
n8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue,
n8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse,
n8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290
BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_left,
BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_right,
BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1
result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1
result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1
result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1
result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_cond,
result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1
result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output);

-- n8_MUX_uxn_opcodes_h_l1331_c7_42b1
n8_MUX_uxn_opcodes_h_l1331_c7_42b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1331_c7_42b1_cond,
n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue,
n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse,
n8_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023
BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_left,
BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_right,
BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef
result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond,
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output);

-- n8_MUX_uxn_opcodes_h_l1334_c7_b2ef
n8_MUX_uxn_opcodes_h_l1334_c7_b2ef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond,
n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue,
n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse,
n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1337_c30_762f
sp_relative_shift_uxn_opcodes_h_l1337_c30_762f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_ins,
sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_x,
sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_y,
sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce
BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_left,
BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_right,
BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_return_output);

-- MUX_uxn_opcodes_h_l1340_c21_7540
MUX_uxn_opcodes_h_l1340_c21_7540 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1340_c21_7540_cond,
MUX_uxn_opcodes_h_l1340_c21_7540_iftrue,
MUX_uxn_opcodes_h_l1340_c21_7540_iffalse,
MUX_uxn_opcodes_h_l1340_c21_7540_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c
BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_left,
BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_right,
BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c
result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c
result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c
result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
 t8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
 n8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output,
 t8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output,
 n8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output,
 t8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output,
 n8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output,
 n8_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output,
 n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output,
 sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_return_output,
 MUX_uxn_opcodes_h_l1340_c21_7540_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1321_c3_5a68 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1320_c3_453d_uxn_opcodes_h_l1320_c3_453d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1325_c3_f076 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1329_c3_7311 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1332_c3_714f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1339_c3_167b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1334_c7_b2ef_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1340_c21_7540_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1340_c21_7540_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1340_c21_7540_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1340_c21_7540_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_0356_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_765b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_0343_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_a467_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1342_DUPLICATE_bf10_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1348_l1315_DUPLICATE_1482_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1329_c3_7311 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1329_c3_7311;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1340_c21_7540_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1332_c3_714f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1332_c3_714f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1321_c3_5a68 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1321_c3_5a68;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1339_c3_167b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1339_c3_167b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1340_c21_7540_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1325_c3_f076 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1325_c3_f076;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1319_c6_a5f2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1331_c11_c290] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_left;
     BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output := BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_0356 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_0356_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_0343 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_0343_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1324_c11_2a30] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_left;
     BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output := BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1327_c11_a578] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_left;
     BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output := BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1337_c30_762f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_ins;
     sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_x;
     sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_return_output := sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_a467 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_a467_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1340_c21_0dce] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_left;
     BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_return_output := BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1342_c11_9c4c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1334_c11_0023] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_left;
     BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output := BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1334_c7_b2ef] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1334_c7_b2ef_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1342_DUPLICATE_bf10 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1342_DUPLICATE_bf10_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_765b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_765b_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c6_a5f2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1324_c11_2a30_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1327_c11_a578_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1331_c11_c290_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1334_c11_0023_return_output;
     VAR_MUX_uxn_opcodes_h_l1340_c21_7540_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1340_c21_0dce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1342_c11_9c4c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_a467_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_a467_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_a467_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_a467_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_a467_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1342_DUPLICATE_bf10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1342_DUPLICATE_bf10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1342_DUPLICATE_bf10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1342_DUPLICATE_bf10_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1342_DUPLICATE_bf10_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_0356_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_0356_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_0356_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_0356_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_0356_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_765b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_765b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_765b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_765b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1331_l1327_l1324_l1319_l1342_DUPLICATE_765b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_0343_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_0343_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_0343_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_0343_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1334_l1331_l1327_l1324_l1319_DUPLICATE_0343_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1334_c7_b2ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1337_c30_762f_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1342_c7_7f0c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1319_c1_46a0] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1327_c7_f738] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1327_c7_f738_cond <= VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_cond;
     t8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue;
     t8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output := t8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;

     -- n8_MUX[uxn_opcodes_h_l1334_c7_b2ef] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond <= VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond;
     n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue;
     n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output := n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1342_c7_7f0c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output;

     -- MUX[uxn_opcodes_h_l1340_c21_7540] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1340_c21_7540_cond <= VAR_MUX_uxn_opcodes_h_l1340_c21_7540_cond;
     MUX_uxn_opcodes_h_l1340_c21_7540_iftrue <= VAR_MUX_uxn_opcodes_h_l1340_c21_7540_iftrue;
     MUX_uxn_opcodes_h_l1340_c21_7540_iffalse <= VAR_MUX_uxn_opcodes_h_l1340_c21_7540_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1340_c21_7540_return_output := MUX_uxn_opcodes_h_l1340_c21_7540_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1334_c7_b2ef] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1342_c7_7f0c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1334_c7_b2ef] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue := VAR_MUX_uxn_opcodes_h_l1340_c21_7540_return_output;
     VAR_printf_uxn_opcodes_h_l1320_c3_453d_uxn_opcodes_h_l1320_c3_453d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1319_c1_46a0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1342_c7_7f0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1334_c7_b2ef] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output := result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1334_c7_b2ef] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1331_c7_42b1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1324_c7_c247] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1324_c7_c247_cond <= VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_cond;
     t8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue;
     t8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output := t8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1334_c7_b2ef] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1334_c7_b2ef] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1331_c7_42b1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1331_c7_42b1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1331_c7_42b1_cond <= VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_cond;
     n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue;
     n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output := n8_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;

     -- printf_uxn_opcodes_h_l1320_c3_453d[uxn_opcodes_h_l1320_c3_453d] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1320_c3_453d_uxn_opcodes_h_l1320_c3_453d_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1320_c3_453d_uxn_opcodes_h_l1320_c3_453d_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1334_c7_b2ef_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1327_c7_f738] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1327_c7_f738] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1331_c7_42b1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1331_c7_42b1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1331_c7_42b1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;

     -- t8_MUX[uxn_opcodes_h_l1319_c2_d110] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1319_c2_d110_cond <= VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_cond;
     t8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue;
     t8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output := t8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1331_c7_42b1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output := result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;

     -- n8_MUX[uxn_opcodes_h_l1327_c7_f738] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1327_c7_f738_cond <= VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_cond;
     n8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue;
     n8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output := n8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1331_c7_42b1_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1324_c7_c247] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1327_c7_f738] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1327_c7_f738] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_return_output := result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1327_c7_f738] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1327_c7_f738] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1324_c7_c247] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;

     -- n8_MUX[uxn_opcodes_h_l1324_c7_c247] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1324_c7_c247_cond <= VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_cond;
     n8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue;
     n8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output := n8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1327_c7_f738_return_output;
     -- n8_MUX[uxn_opcodes_h_l1319_c2_d110] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1319_c2_d110_cond <= VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_cond;
     n8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue;
     n8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output := n8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1319_c2_d110] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1324_c7_c247] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1324_c7_c247] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1324_c7_c247] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_return_output := result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1319_c2_d110] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1324_c7_c247] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1324_c7_c247_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1319_c2_d110] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1319_c2_d110] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_return_output := result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1319_c2_d110] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1319_c2_d110] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1348_l1315_DUPLICATE_1482 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1348_l1315_DUPLICATE_1482_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c2_d110_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c2_d110_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1348_l1315_DUPLICATE_1482_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1348_l1315_DUPLICATE_1482_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
