-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity and_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_bacf6a1d;
architecture arch of and_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l877_c6_1df3]
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l877_c1_3e56]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l877_c2_b935]
signal n8_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l877_c2_b935]
signal t8_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l877_c2_b935]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l877_c2_b935]
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c2_b935]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l877_c2_b935]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l877_c2_b935]
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l877_c2_b935]
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l878_c3_5f4f[uxn_opcodes_h_l878_c3_5f4f]
signal printf_uxn_opcodes_h_l878_c3_5f4f_uxn_opcodes_h_l878_c3_5f4f_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l882_c11_6b02]
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l882_c7_b288]
signal n8_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l882_c7_b288]
signal t8_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l882_c7_b288]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l882_c7_b288]
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l882_c7_b288]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l882_c7_b288]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l882_c7_b288]
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l882_c7_b288]
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l885_c11_e969]
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l885_c7_ef5b]
signal n8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l885_c7_ef5b]
signal t8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l885_c7_ef5b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l885_c7_ef5b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l885_c7_ef5b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l885_c7_ef5b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l885_c7_ef5b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l885_c7_ef5b]
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l888_c11_3d18]
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l888_c7_cb2f]
signal n8_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l888_c7_cb2f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l888_c7_cb2f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l888_c7_cb2f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l888_c7_cb2f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l888_c7_cb2f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l888_c7_cb2f]
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l891_c30_63fb]
signal sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l894_c21_d1c8]
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l896_c11_cf77]
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l896_c7_a36f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l896_c7_a36f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l896_c7_a36f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4e73( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3
BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_left,
BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_right,
BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_return_output);

-- n8_MUX_uxn_opcodes_h_l877_c2_b935
n8_MUX_uxn_opcodes_h_l877_c2_b935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l877_c2_b935_cond,
n8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue,
n8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse,
n8_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

-- t8_MUX_uxn_opcodes_h_l877_c2_b935
t8_MUX_uxn_opcodes_h_l877_c2_b935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l877_c2_b935_cond,
t8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue,
t8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse,
t8_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935
result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_cond,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

-- printf_uxn_opcodes_h_l878_c3_5f4f_uxn_opcodes_h_l878_c3_5f4f
printf_uxn_opcodes_h_l878_c3_5f4f_uxn_opcodes_h_l878_c3_5f4f : entity work.printf_uxn_opcodes_h_l878_c3_5f4f_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l878_c3_5f4f_uxn_opcodes_h_l878_c3_5f4f_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02
BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_left,
BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_right,
BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output);

-- n8_MUX_uxn_opcodes_h_l882_c7_b288
n8_MUX_uxn_opcodes_h_l882_c7_b288 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l882_c7_b288_cond,
n8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue,
n8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse,
n8_MUX_uxn_opcodes_h_l882_c7_b288_return_output);

-- t8_MUX_uxn_opcodes_h_l882_c7_b288
t8_MUX_uxn_opcodes_h_l882_c7_b288 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l882_c7_b288_cond,
t8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue,
t8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse,
t8_MUX_uxn_opcodes_h_l882_c7_b288_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288
result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_cond,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969
BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_left,
BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_right,
BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output);

-- n8_MUX_uxn_opcodes_h_l885_c7_ef5b
n8_MUX_uxn_opcodes_h_l885_c7_ef5b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond,
n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue,
n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse,
n8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output);

-- t8_MUX_uxn_opcodes_h_l885_c7_ef5b
t8_MUX_uxn_opcodes_h_l885_c7_ef5b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond,
t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue,
t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse,
t8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b
result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_cond,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18
BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_left,
BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_right,
BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output);

-- n8_MUX_uxn_opcodes_h_l888_c7_cb2f
n8_MUX_uxn_opcodes_h_l888_c7_cb2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l888_c7_cb2f_cond,
n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue,
n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse,
n8_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f
result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_cond,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l891_c30_63fb
sp_relative_shift_uxn_opcodes_h_l891_c30_63fb : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_ins,
sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_x,
sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_y,
sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8
BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_left,
BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_right,
BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77
BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_left,
BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_right,
BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_return_output,
 n8_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
 t8_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output,
 n8_MUX_uxn_opcodes_h_l882_c7_b288_return_output,
 t8_MUX_uxn_opcodes_h_l882_c7_b288_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output,
 n8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output,
 t8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output,
 n8_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output,
 sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_return_output,
 BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_6d08 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l878_c3_5f4f_uxn_opcodes_h_l878_c3_5f4f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_87b0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_c09a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_c0ff_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_d382_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_191c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_bcea_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l885_l888_l882_l896_DUPLICATE_bbcc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_7c20_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l873_l902_DUPLICATE_db7d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_87b0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_87b0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_6d08 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_6d08;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_c09a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_c09a;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l896_c11_cf77] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_left;
     BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output := BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_191c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_191c_return_output := result.sp_relative_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l894_c21_d1c8] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_left;
     BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_return_output := BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l891_c30_63fb] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_ins;
     sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_x <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_x;
     sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_y <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_return_output := sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_d382 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_d382_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_c0ff LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_c0ff_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_bcea LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_bcea_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l882_c11_6b02] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_left;
     BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output := BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l888_c11_3d18] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_left;
     BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output := BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l885_c11_e969] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_left;
     BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output := BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l877_c6_1df3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_left;
     BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output := BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l885_l888_l882_l896_DUPLICATE_bbcc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l885_l888_l882_l896_DUPLICATE_bbcc_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_7c20 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_7c20_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_d1c8_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_1df3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_6b02_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_e969_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3d18_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_cf77_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_191c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_191c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_191c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_191c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l885_l888_l882_l896_DUPLICATE_bbcc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l885_l888_l882_l896_DUPLICATE_bbcc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l885_l888_l882_l896_DUPLICATE_bbcc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l885_l888_l882_l896_DUPLICATE_bbcc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_d382_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_d382_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_d382_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_d382_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_c0ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_c0ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_c0ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l885_l877_l882_l896_DUPLICATE_c0ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_7c20_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_7c20_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_bcea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_bcea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_bcea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l885_l877_l888_l882_DUPLICATE_bcea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_63fb_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l888_c7_cb2f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output := result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;

     -- t8_MUX[uxn_opcodes_h_l885_c7_ef5b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond;
     t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue;
     t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output := t8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l896_c7_a36f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l877_c1_3e56] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l896_c7_a36f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l888_c7_cb2f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l896_c7_a36f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_return_output;

     -- n8_MUX[uxn_opcodes_h_l888_c7_cb2f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l888_c7_cb2f_cond <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_cond;
     n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue;
     n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output := n8_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l888_c7_cb2f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l878_c3_5f4f_uxn_opcodes_h_l878_c3_5f4f_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_3e56_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_a36f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_a36f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_a36f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse := VAR_t8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l885_c7_ef5b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;

     -- n8_MUX[uxn_opcodes_h_l885_c7_ef5b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_cond;
     n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue;
     n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output := n8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l885_c7_ef5b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l888_c7_cb2f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;

     -- t8_MUX[uxn_opcodes_h_l882_c7_b288] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l882_c7_b288_cond <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_cond;
     t8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue;
     t8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_return_output := t8_MUX_uxn_opcodes_h_l882_c7_b288_return_output;

     -- printf_uxn_opcodes_h_l878_c3_5f4f[uxn_opcodes_h_l878_c3_5f4f] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l878_c3_5f4f_uxn_opcodes_h_l878_c3_5f4f_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l878_c3_5f4f_uxn_opcodes_h_l878_c3_5f4f_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l885_c7_ef5b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output := result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l888_c7_cb2f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l888_c7_cb2f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse := VAR_n8_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_cb2f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse := VAR_t8_MUX_uxn_opcodes_h_l882_c7_b288_return_output;
     -- t8_MUX[uxn_opcodes_h_l877_c2_b935] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l877_c2_b935_cond <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_cond;
     t8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue;
     t8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_return_output := t8_MUX_uxn_opcodes_h_l877_c2_b935_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l885_c7_ef5b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l882_c7_b288] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l885_c7_ef5b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;

     -- n8_MUX[uxn_opcodes_h_l882_c7_b288] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l882_c7_b288_cond <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_cond;
     n8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_iftrue;
     n8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_return_output := n8_MUX_uxn_opcodes_h_l882_c7_b288_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l882_c7_b288] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l885_c7_ef5b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l882_c7_b288] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_cond;
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_return_output := result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse := VAR_n8_MUX_uxn_opcodes_h_l882_c7_b288_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_ef5b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_b288_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_b288_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l877_c2_b935_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l882_c7_b288] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l877_c2_b935] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l877_c2_b935] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_cond;
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_return_output := result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_return_output;

     -- n8_MUX[uxn_opcodes_h_l877_c2_b935] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l877_c2_b935_cond <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_cond;
     n8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_iftrue;
     n8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_return_output := n8_MUX_uxn_opcodes_h_l877_c2_b935_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l877_c2_b935] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l882_c7_b288] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l882_c7_b288] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l877_c2_b935_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_b288_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_b288_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_b288_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c2_b935] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l877_c2_b935] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l877_c2_b935] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l873_l902_DUPLICATE_db7d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l873_l902_DUPLICATE_db7d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4e73(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_b935_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_b935_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l873_l902_DUPLICATE_db7d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l873_l902_DUPLICATE_db7d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
