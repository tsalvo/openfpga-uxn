-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 37
entity dup_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_6be78140;
architecture arch of dup_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2608_c6_fddc]
signal BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2608_c1_7d78]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2608_c2_95f2]
signal t8_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2608_c2_95f2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2608_c2_95f2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2608_c2_95f2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2608_c2_95f2]
signal result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2608_c2_95f2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2608_c2_95f2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(0 downto 0);

-- printf_uxn_opcodes_h_l2609_c3_0e00[uxn_opcodes_h_l2609_c3_0e00]
signal printf_uxn_opcodes_h_l2609_c3_0e00_uxn_opcodes_h_l2609_c3_0e00_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2613_c11_2efd]
signal BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2613_c7_77fa]
signal t8_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2613_c7_77fa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2613_c7_77fa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2613_c7_77fa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2613_c7_77fa]
signal result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2613_c7_77fa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2613_c7_77fa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2616_c11_8203]
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2616_c7_e164]
signal t8_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2616_c7_e164]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2616_c7_e164]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2616_c7_e164]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2616_c7_e164]
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2616_c7_e164]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2616_c7_e164]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2619_c30_341e]
signal sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2624_c11_e5f4]
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2624_c7_9f75]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2624_c7_9f75]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2624_c7_9f75]
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2624_c7_9f75]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2624_c7_9f75]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2629_c11_ae44]
signal BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2629_c7_995b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2629_c7_995b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c551( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc
BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_left,
BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_right,
BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_return_output);

-- t8_MUX_uxn_opcodes_h_l2608_c2_95f2
t8_MUX_uxn_opcodes_h_l2608_c2_95f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2608_c2_95f2_cond,
t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue,
t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse,
t8_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2
result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2
result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2
result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2
result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2
result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output);

-- printf_uxn_opcodes_h_l2609_c3_0e00_uxn_opcodes_h_l2609_c3_0e00
printf_uxn_opcodes_h_l2609_c3_0e00_uxn_opcodes_h_l2609_c3_0e00 : entity work.printf_uxn_opcodes_h_l2609_c3_0e00_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2609_c3_0e00_uxn_opcodes_h_l2609_c3_0e00_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd
BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_left,
BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_right,
BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output);

-- t8_MUX_uxn_opcodes_h_l2613_c7_77fa
t8_MUX_uxn_opcodes_h_l2613_c7_77fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2613_c7_77fa_cond,
t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue,
t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse,
t8_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa
result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa
result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa
result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_cond,
result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa
result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa
result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203
BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_left,
BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_right,
BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output);

-- t8_MUX_uxn_opcodes_h_l2616_c7_e164
t8_MUX_uxn_opcodes_h_l2616_c7_e164 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2616_c7_e164_cond,
t8_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue,
t8_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse,
t8_MUX_uxn_opcodes_h_l2616_c7_e164_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_cond,
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2619_c30_341e
sp_relative_shift_uxn_opcodes_h_l2619_c30_341e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_ins,
sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_x,
sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_y,
sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_left,
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_right,
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_cond,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44
BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_left,
BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_right,
BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b
result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b
result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_return_output,
 t8_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output,
 t8_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output,
 t8_MUX_uxn_opcodes_h_l2616_c7_e164_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output,
 sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2610_c3_b9a3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2609_c3_0e00_uxn_opcodes_h_l2609_c3_0e00_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2614_c3_937f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_cc4a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_0c0f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2624_c7_9f75_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2608_DUPLICATE_038e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2613_l2616_l2608_DUPLICATE_a90e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_5908_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_1c5f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2616_DUPLICATE_914e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2634_l2604_DUPLICATE_35c1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2610_c3_b9a3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2610_c3_b9a3;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_0c0f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2626_c3_0c0f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_cc4a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2621_c3_cc4a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2614_c3_937f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2614_c3_937f;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2608_DUPLICATE_038e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2608_DUPLICATE_038e_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2629_c11_ae44] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_left;
     BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_return_output := BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2624_c11_e5f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_1c5f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_1c5f_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2616_c11_8203] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_left;
     BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output := BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2619_c30_341e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_ins;
     sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_x;
     sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_return_output := sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2624_c7_9f75] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2624_c7_9f75_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_5908 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_5908_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2608_c6_fddc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_left;
     BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output := BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2613_c11_2efd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2613_l2616_l2608_DUPLICATE_a90e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2613_l2616_l2608_DUPLICATE_a90e_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2616_DUPLICATE_914e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2616_DUPLICATE_914e_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2608_c6_fddc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2613_c11_2efd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c11_8203_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_e5f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2629_c11_ae44_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2613_l2616_l2608_DUPLICATE_a90e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2613_l2616_l2608_DUPLICATE_a90e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2613_l2616_l2608_DUPLICATE_a90e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2616_DUPLICATE_914e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2616_DUPLICATE_914e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2616_DUPLICATE_914e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2616_DUPLICATE_914e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_1c5f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_1c5f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_1c5f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2608_DUPLICATE_038e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2608_DUPLICATE_038e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2608_DUPLICATE_038e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2624_l2613_l2629_l2608_DUPLICATE_038e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_5908_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_5908_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2624_l2613_l2608_DUPLICATE_5908_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2624_c7_9f75_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2619_c30_341e_return_output;
     -- t8_MUX[uxn_opcodes_h_l2616_c7_e164] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2616_c7_e164_cond <= VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_cond;
     t8_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue;
     t8_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_return_output := t8_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2616_c7_e164] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2624_c7_9f75] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2629_c7_995b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2608_c1_7d78] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2624_c7_9f75] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2629_c7_995b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2624_c7_9f75] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output := result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2609_c3_0e00_uxn_opcodes_h_l2609_c3_0e00_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2608_c1_7d78_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2629_c7_995b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2629_c7_995b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2616_c7_e164] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_return_output := result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;

     -- t8_MUX[uxn_opcodes_h_l2613_c7_77fa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2613_c7_77fa_cond <= VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_cond;
     t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue;
     t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output := t8_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2613_c7_77fa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;

     -- printf_uxn_opcodes_h_l2609_c3_0e00[uxn_opcodes_h_l2609_c3_0e00] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2609_c3_0e00_uxn_opcodes_h_l2609_c3_0e00_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2609_c3_0e00_uxn_opcodes_h_l2609_c3_0e00_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2616_c7_e164] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2624_c7_9f75] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2616_c7_e164] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2624_c7_9f75] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_9f75_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2616_c7_e164] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2608_c2_95f2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2613_c7_77fa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2616_c7_e164] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;

     -- t8_MUX[uxn_opcodes_h_l2608_c2_95f2] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2608_c2_95f2_cond <= VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_cond;
     t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue;
     t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output := t8_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2613_c7_77fa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output := result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2613_c7_77fa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c7_e164_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2613_c7_77fa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2608_c2_95f2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2608_c2_95f2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2613_c7_77fa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2608_c2_95f2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2613_c7_77fa_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2608_c2_95f2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2608_c2_95f2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2634_l2604_DUPLICATE_35c1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2634_l2604_DUPLICATE_35c1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c551(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2608_c2_95f2_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2634_l2604_DUPLICATE_35c1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c551_uxn_opcodes_h_l2634_l2604_DUPLICATE_35c1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
