-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity neq_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_6d7675a8;
architecture arch of neq_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1314_c6_a19b]
signal BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1314_c1_0672]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1314_c2_e6bf]
signal n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1314_c2_e6bf]
signal t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1314_c2_e6bf]
signal result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1314_c2_e6bf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1314_c2_e6bf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1314_c2_e6bf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1314_c2_e6bf]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1314_c2_e6bf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(3 downto 0);

-- printf_uxn_opcodes_h_l1315_c3_5bfc[uxn_opcodes_h_l1315_c3_5bfc]
signal printf_uxn_opcodes_h_l1315_c3_5bfc_uxn_opcodes_h_l1315_c3_5bfc_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1319_c11_1c51]
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1319_c7_f274]
signal n8_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1319_c7_f274]
signal t8_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1319_c7_f274]
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1319_c7_f274]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1319_c7_f274]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1319_c7_f274]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1319_c7_f274]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1319_c7_f274]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1322_c11_decb]
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1322_c7_d1f4]
signal n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1322_c7_d1f4]
signal t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1322_c7_d1f4]
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1322_c7_d1f4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1322_c7_d1f4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1322_c7_d1f4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1322_c7_d1f4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1322_c7_d1f4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1326_c11_e8a6]
signal BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1326_c7_91e2]
signal n8_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1326_c7_91e2]
signal result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1326_c7_91e2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1326_c7_91e2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1326_c7_91e2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1326_c7_91e2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1326_c7_91e2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1329_c11_74de]
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1329_c7_f741]
signal n8_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1329_c7_f741]
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1329_c7_f741]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1329_c7_f741]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1329_c7_f741]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1329_c7_f741]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1329_c7_f741]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1332_c30_4507]
signal sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1335_c21_2d65]
signal BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1335_c21_f37c]
signal MUX_uxn_opcodes_h_l1335_c21_f37c_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1335_c21_f37c_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1335_c21_f37c_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1335_c21_f37c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1337_c11_ba08]
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1337_c7_118e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1337_c7_118e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1337_c7_118e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_25e8( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b
BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_left,
BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_right,
BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_return_output);

-- n8_MUX_uxn_opcodes_h_l1314_c2_e6bf
n8_MUX_uxn_opcodes_h_l1314_c2_e6bf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond,
n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue,
n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse,
n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

-- t8_MUX_uxn_opcodes_h_l1314_c2_e6bf
t8_MUX_uxn_opcodes_h_l1314_c2_e6bf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond,
t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue,
t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse,
t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond,
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

-- printf_uxn_opcodes_h_l1315_c3_5bfc_uxn_opcodes_h_l1315_c3_5bfc
printf_uxn_opcodes_h_l1315_c3_5bfc_uxn_opcodes_h_l1315_c3_5bfc : entity work.printf_uxn_opcodes_h_l1315_c3_5bfc_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1315_c3_5bfc_uxn_opcodes_h_l1315_c3_5bfc_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51
BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_left,
BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_right,
BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output);

-- n8_MUX_uxn_opcodes_h_l1319_c7_f274
n8_MUX_uxn_opcodes_h_l1319_c7_f274 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1319_c7_f274_cond,
n8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue,
n8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse,
n8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output);

-- t8_MUX_uxn_opcodes_h_l1319_c7_f274
t8_MUX_uxn_opcodes_h_l1319_c7_f274 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1319_c7_f274_cond,
t8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue,
t8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse,
t8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_cond,
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_left,
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_right,
BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output);

-- n8_MUX_uxn_opcodes_h_l1322_c7_d1f4
n8_MUX_uxn_opcodes_h_l1322_c7_d1f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond,
n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue,
n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse,
n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output);

-- t8_MUX_uxn_opcodes_h_l1322_c7_d1f4
t8_MUX_uxn_opcodes_h_l1322_c7_d1f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond,
t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue,
t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse,
t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6
BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_left,
BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_right,
BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output);

-- n8_MUX_uxn_opcodes_h_l1326_c7_91e2
n8_MUX_uxn_opcodes_h_l1326_c7_91e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1326_c7_91e2_cond,
n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue,
n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse,
n8_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_left,
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_right,
BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output);

-- n8_MUX_uxn_opcodes_h_l1329_c7_f741
n8_MUX_uxn_opcodes_h_l1329_c7_f741 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1329_c7_f741_cond,
n8_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue,
n8_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse,
n8_MUX_uxn_opcodes_h_l1329_c7_f741_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_cond,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1332_c30_4507
sp_relative_shift_uxn_opcodes_h_l1332_c30_4507 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_ins,
sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_x,
sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_y,
sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65
BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_left,
BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_right,
BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_return_output);

-- MUX_uxn_opcodes_h_l1335_c21_f37c
MUX_uxn_opcodes_h_l1335_c21_f37c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1335_c21_f37c_cond,
MUX_uxn_opcodes_h_l1335_c21_f37c_iftrue,
MUX_uxn_opcodes_h_l1335_c21_f37c_iffalse,
MUX_uxn_opcodes_h_l1335_c21_f37c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_left,
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_right,
BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_return_output,
 n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
 t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output,
 n8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output,
 t8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output,
 n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output,
 t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output,
 n8_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output,
 n8_MUX_uxn_opcodes_h_l1329_c7_f741_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_return_output,
 sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_return_output,
 MUX_uxn_opcodes_h_l1335_c21_f37c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1316_c3_8d62 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1315_c3_5bfc_uxn_opcodes_h_l1315_c3_5bfc_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1320_c3_8fbe : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1324_c3_c013 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_89ce : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1334_c3_0b0f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1329_c7_f741_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_c854_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_b933_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_3590_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_875d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1337_l1329_l1326_l1322_l1319_DUPLICATE_3e56_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1343_l1310_DUPLICATE_db9e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1316_c3_8d62 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1316_c3_8d62;
     VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1334_c3_0b0f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1334_c3_0b0f;
     VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1320_c3_8fbe := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1320_c3_8fbe;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1324_c3_c013 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1324_c3_c013;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_89ce := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1327_c3_89ce;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_3590 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_3590_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1337_l1329_l1326_l1322_l1319_DUPLICATE_3e56 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1337_l1329_l1326_l1322_l1319_DUPLICATE_3e56_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1326_c11_e8a6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_b933 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_b933_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_c854 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_c854_return_output := result.u8_value;

     -- sp_relative_shift[uxn_opcodes_h_l1332_c30_4507] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_ins;
     sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_x;
     sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_return_output := sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1329_c7_f741] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1329_c7_f741_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1337_c11_ba08] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_left;
     BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output := BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1322_c11_decb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_left;
     BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output := BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1335_c21_2d65] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_left;
     BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_return_output := BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1314_c6_a19b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_875d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_875d_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1329_c11_74de] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_left;
     BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output := BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1319_c11_1c51] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_left;
     BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output := BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1314_c6_a19b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1319_c11_1c51_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1322_c11_decb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1326_c11_e8a6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1329_c11_74de_return_output;
     VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1335_c21_2d65_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1337_c11_ba08_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_b933_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_b933_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_b933_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_b933_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_b933_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1337_l1329_l1326_l1322_l1319_DUPLICATE_3e56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1337_l1329_l1326_l1322_l1319_DUPLICATE_3e56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1337_l1329_l1326_l1322_l1319_DUPLICATE_3e56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1337_l1329_l1326_l1322_l1319_DUPLICATE_3e56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1337_l1329_l1326_l1322_l1319_DUPLICATE_3e56_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_875d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_875d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_875d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_875d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_875d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_3590_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_3590_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_3590_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_3590_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1337_l1326_l1322_l1319_l1314_DUPLICATE_3590_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_c854_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_c854_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_c854_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_c854_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1329_l1326_l1322_l1319_l1314_DUPLICATE_c854_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1329_c7_f741_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1332_c30_4507_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1329_c7_f741] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1337_c7_118e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_return_output;

     -- t8_MUX[uxn_opcodes_h_l1322_c7_d1f4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond;
     t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue;
     t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output := t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1329_c7_f741] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;

     -- n8_MUX[uxn_opcodes_h_l1329_c7_f741] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1329_c7_f741_cond <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_cond;
     n8_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue;
     n8_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_return_output := n8_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1337_c7_118e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_return_output;

     -- MUX[uxn_opcodes_h_l1335_c21_f37c] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1335_c21_f37c_cond <= VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_cond;
     MUX_uxn_opcodes_h_l1335_c21_f37c_iftrue <= VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_iftrue;
     MUX_uxn_opcodes_h_l1335_c21_f37c_iffalse <= VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_return_output := MUX_uxn_opcodes_h_l1335_c21_f37c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1314_c1_0672] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1337_c7_118e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue := VAR_MUX_uxn_opcodes_h_l1335_c21_f37c_return_output;
     VAR_printf_uxn_opcodes_h_l1315_c3_5bfc_uxn_opcodes_h_l1315_c3_5bfc_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1314_c1_0672_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1337_c7_118e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1337_c7_118e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1337_c7_118e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1329_c7_f741] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1326_c7_91e2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1329_c7_f741] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1329_c7_f741] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;

     -- t8_MUX[uxn_opcodes_h_l1319_c7_f274] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1319_c7_f274_cond <= VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_cond;
     t8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue;
     t8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output := t8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1326_c7_91e2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;

     -- printf_uxn_opcodes_h_l1315_c3_5bfc[uxn_opcodes_h_l1315_c3_5bfc] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1315_c3_5bfc_uxn_opcodes_h_l1315_c3_5bfc_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1315_c3_5bfc_uxn_opcodes_h_l1315_c3_5bfc_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_u8_value_MUX[uxn_opcodes_h_l1329_c7_f741] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_return_output := result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;

     -- n8_MUX[uxn_opcodes_h_l1326_c7_91e2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1326_c7_91e2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_cond;
     n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue;
     n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output := n8_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1329_c7_f741_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1326_c7_91e2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1326_c7_91e2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1322_c7_d1f4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1326_c7_91e2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;

     -- t8_MUX[uxn_opcodes_h_l1314_c2_e6bf] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond <= VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond;
     t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue;
     t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output := t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1326_c7_91e2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1322_c7_d1f4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1322_c7_d1f4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond;
     n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue;
     n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output := n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1326_c7_91e2_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1322_c7_d1f4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1322_c7_d1f4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1319_c7_f274] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1319_c7_f274_cond <= VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_cond;
     n8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue;
     n8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output := n8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1322_c7_d1f4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1319_c7_f274] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1322_c7_d1f4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1319_c7_f274] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1322_c7_d1f4_return_output;
     -- n8_MUX[uxn_opcodes_h_l1314_c2_e6bf] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond <= VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond;
     n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue;
     n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output := n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1319_c7_f274] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1319_c7_f274] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_return_output := result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1314_c2_e6bf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1319_c7_f274] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1319_c7_f274] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1314_c2_e6bf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1319_c7_f274_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1314_c2_e6bf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1314_c2_e6bf] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1314_c2_e6bf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output := result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1314_c2_e6bf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1343_l1310_DUPLICATE_db9e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1343_l1310_DUPLICATE_db9e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_25e8(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1314_c2_e6bf_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1343_l1310_DUPLICATE_db9e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_25e8_uxn_opcodes_h_l1343_l1310_DUPLICATE_db9e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
