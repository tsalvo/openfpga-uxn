-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity jmp2_0CLK_355c9936 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jmp2_0CLK_355c9936;
architecture arch of jmp2_0CLK_355c9936 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l652_c6_4b1a]
signal BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l652_c2_885b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l652_c2_885b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l652_c2_885b]
signal result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l652_c2_885b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l652_c2_885b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l652_c2_885b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l652_c2_885b]
signal t16_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l657_c11_016d]
signal BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l657_c7_63c9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l657_c7_63c9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l657_c7_63c9]
signal result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l657_c7_63c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l657_c7_63c9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l657_c7_63c9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l657_c7_63c9]
signal t16_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l660_c11_10dd]
signal BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l660_c7_1479]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l660_c7_1479]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l660_c7_1479]
signal result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l660_c7_1479]
signal result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l660_c7_1479]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l660_c7_1479]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l660_c7_1479]
signal t16_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l662_c3_c19b]
signal CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l665_c11_635b]
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l665_c7_f085]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l665_c7_f085]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l665_c7_f085]
signal result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l665_c7_f085]
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l665_c7_f085]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l665_c7_f085]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l665_c7_f085]
signal t16_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l668_c11_163b]
signal BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l668_c7_b910]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l668_c7_b910]
signal result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l668_c7_b910]
signal result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l668_c7_b910]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l668_c7_b910]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l668_c7_b910]
signal t16_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l669_c3_de1f]
signal BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l671_c30_8964]
signal sp_relative_shift_uxn_opcodes_h_l671_c30_8964_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l671_c30_8964_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l671_c30_8964_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l671_c30_8964_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l675_c11_ec62]
signal BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l675_c7_da6a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l675_c7_da6a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l675_c7_da6a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a
BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_left,
BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_right,
BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b
result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_cond,
result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output);

-- t16_MUX_uxn_opcodes_h_l652_c2_885b
t16_MUX_uxn_opcodes_h_l652_c2_885b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l652_c2_885b_cond,
t16_MUX_uxn_opcodes_h_l652_c2_885b_iftrue,
t16_MUX_uxn_opcodes_h_l652_c2_885b_iffalse,
t16_MUX_uxn_opcodes_h_l652_c2_885b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d
BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_left,
BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_right,
BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9
result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_cond,
result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output);

-- t16_MUX_uxn_opcodes_h_l657_c7_63c9
t16_MUX_uxn_opcodes_h_l657_c7_63c9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l657_c7_63c9_cond,
t16_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue,
t16_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse,
t16_MUX_uxn_opcodes_h_l657_c7_63c9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd
BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_left,
BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_right,
BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479
result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_cond,
result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output);

-- t16_MUX_uxn_opcodes_h_l660_c7_1479
t16_MUX_uxn_opcodes_h_l660_c7_1479 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l660_c7_1479_cond,
t16_MUX_uxn_opcodes_h_l660_c7_1479_iftrue,
t16_MUX_uxn_opcodes_h_l660_c7_1479_iffalse,
t16_MUX_uxn_opcodes_h_l660_c7_1479_return_output);

-- CONST_SL_8_uxn_opcodes_h_l662_c3_c19b
CONST_SL_8_uxn_opcodes_h_l662_c3_c19b : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_x,
CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b
BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_left,
BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_right,
BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085
result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_cond,
result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output);

-- t16_MUX_uxn_opcodes_h_l665_c7_f085
t16_MUX_uxn_opcodes_h_l665_c7_f085 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l665_c7_f085_cond,
t16_MUX_uxn_opcodes_h_l665_c7_f085_iftrue,
t16_MUX_uxn_opcodes_h_l665_c7_f085_iffalse,
t16_MUX_uxn_opcodes_h_l665_c7_f085_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b
BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_left,
BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_right,
BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910
result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_cond,
result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output);

-- t16_MUX_uxn_opcodes_h_l668_c7_b910
t16_MUX_uxn_opcodes_h_l668_c7_b910 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l668_c7_b910_cond,
t16_MUX_uxn_opcodes_h_l668_c7_b910_iftrue,
t16_MUX_uxn_opcodes_h_l668_c7_b910_iffalse,
t16_MUX_uxn_opcodes_h_l668_c7_b910_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f
BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_left,
BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_right,
BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l671_c30_8964
sp_relative_shift_uxn_opcodes_h_l671_c30_8964 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l671_c30_8964_ins,
sp_relative_shift_uxn_opcodes_h_l671_c30_8964_x,
sp_relative_shift_uxn_opcodes_h_l671_c30_8964_y,
sp_relative_shift_uxn_opcodes_h_l671_c30_8964_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62
BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_left,
BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_right,
BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
 t16_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output,
 t16_MUX_uxn_opcodes_h_l657_c7_63c9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output,
 t16_MUX_uxn_opcodes_h_l660_c7_1479_return_output,
 CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output,
 t16_MUX_uxn_opcodes_h_l665_c7_f085_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output,
 t16_MUX_uxn_opcodes_h_l668_c7_b910_return_output,
 BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_return_output,
 sp_relative_shift_uxn_opcodes_h_l671_c30_8964_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l654_c3_2a8b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_ed1c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l663_c3_c017 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l666_c3_edde : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l665_c7_f085_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_f56b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_76f5_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_07c3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_47d5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l668_l657_l675_DUPLICATE_45dd_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l661_l669_DUPLICATE_fb26_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l681_l648_DUPLICATE_1d01_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l663_c3_c017 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l663_c3_c017;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l666_c3_edde := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l666_c3_edde;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_ed1c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l658_c3_ed1c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l654_c3_2a8b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l654_c3_2a8b;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_y := resize(to_signed(-2, 3), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l657_c11_016d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_left;
     BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output := BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_f56b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_f56b_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l668_c11_163b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_left;
     BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output := BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l652_c6_4b1a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_left;
     BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output := BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l671_c30_8964] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l671_c30_8964_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_ins;
     sp_relative_shift_uxn_opcodes_h_l671_c30_8964_x <= VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_x;
     sp_relative_shift_uxn_opcodes_h_l671_c30_8964_y <= VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_return_output := sp_relative_shift_uxn_opcodes_h_l671_c30_8964_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l675_c11_ec62] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_left;
     BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output := BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_07c3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_07c3_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l665_c11_635b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_left;
     BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output := BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l661_l669_DUPLICATE_fb26 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l661_l669_DUPLICATE_fb26_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l660_c11_10dd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_left;
     BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output := BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l668_l657_l675_DUPLICATE_45dd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l668_l657_l675_DUPLICATE_45dd_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_76f5 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_76f5_return_output := result.u16_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l665_c7_f085] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l665_c7_f085_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_47d5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_47d5_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l652_c6_4b1a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l657_c11_016d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l660_c11_10dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_635b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l668_c11_163b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l675_c11_ec62_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l661_l669_DUPLICATE_fb26_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l661_l669_DUPLICATE_fb26_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_07c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_07c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_07c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_07c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_07c3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_76f5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_76f5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_76f5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_76f5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l660_l665_l652_l668_l657_DUPLICATE_76f5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l668_l657_l675_DUPLICATE_45dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l668_l657_l675_DUPLICATE_45dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l668_l657_l675_DUPLICATE_45dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l668_l657_l675_DUPLICATE_45dd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l660_l665_l668_l657_l675_DUPLICATE_45dd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_f56b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_f56b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_f56b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_f56b_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_f56b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_47d5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_47d5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_47d5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_47d5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l660_l665_l652_l657_l675_DUPLICATE_47d5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l665_c7_f085_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l671_c30_8964_return_output;
     -- BIN_OP_OR[uxn_opcodes_h_l669_c3_de1f] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_left;
     BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_return_output := BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l662_c3_c19b] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_x <= VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_return_output := CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l665_c7_f085] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l668_c7_b910] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l675_c7_da6a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l675_c7_da6a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l675_c7_da6a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l669_c3_de1f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l662_c3_c19b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l675_c7_da6a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l675_c7_da6a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l675_c7_da6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l665_c7_f085_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l660_c7_1479] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_return_output;

     -- t16_MUX[uxn_opcodes_h_l668_c7_b910] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l668_c7_b910_cond <= VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_cond;
     t16_MUX_uxn_opcodes_h_l668_c7_b910_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_iftrue;
     t16_MUX_uxn_opcodes_h_l668_c7_b910_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_return_output := t16_MUX_uxn_opcodes_h_l668_c7_b910_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l668_c7_b910] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_cond;
     result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_return_output := result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l668_c7_b910] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l668_c7_b910] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l668_c7_b910] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l665_c7_f085] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l668_c7_b910_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l668_c7_b910_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l668_c7_b910_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l660_c7_1479_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l668_c7_b910_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_iffalse := VAR_t16_MUX_uxn_opcodes_h_l668_c7_b910_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l657_c7_63c9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l665_c7_f085] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output;

     -- t16_MUX[uxn_opcodes_h_l665_c7_f085] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l665_c7_f085_cond <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_cond;
     t16_MUX_uxn_opcodes_h_l665_c7_f085_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_iftrue;
     t16_MUX_uxn_opcodes_h_l665_c7_f085_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_return_output := t16_MUX_uxn_opcodes_h_l665_c7_f085_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l665_c7_f085] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l665_c7_f085] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_cond;
     result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_return_output := result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l665_c7_f085] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l660_c7_1479] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_f085_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_f085_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l665_c7_f085_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_f085_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_iffalse := VAR_t16_MUX_uxn_opcodes_h_l665_c7_f085_return_output;
     -- t16_MUX[uxn_opcodes_h_l660_c7_1479] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l660_c7_1479_cond <= VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_cond;
     t16_MUX_uxn_opcodes_h_l660_c7_1479_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_iftrue;
     t16_MUX_uxn_opcodes_h_l660_c7_1479_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_return_output := t16_MUX_uxn_opcodes_h_l660_c7_1479_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l660_c7_1479] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l660_c7_1479] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_cond;
     result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_return_output := result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l660_c7_1479] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l660_c7_1479] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l657_c7_63c9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l652_c2_885b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l660_c7_1479_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l660_c7_1479_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l660_c7_1479_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l660_c7_1479_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse := VAR_t16_MUX_uxn_opcodes_h_l660_c7_1479_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l657_c7_63c9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_return_output := result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l652_c2_885b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l657_c7_63c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l657_c7_63c9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;

     -- t16_MUX[uxn_opcodes_h_l657_c7_63c9] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l657_c7_63c9_cond <= VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_cond;
     t16_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue;
     t16_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_return_output := t16_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l657_c7_63c9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_iffalse := VAR_t16_MUX_uxn_opcodes_h_l657_c7_63c9_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l652_c2_885b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l652_c2_885b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_return_output;

     -- t16_MUX[uxn_opcodes_h_l652_c2_885b] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l652_c2_885b_cond <= VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_cond;
     t16_MUX_uxn_opcodes_h_l652_c2_885b_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_iftrue;
     t16_MUX_uxn_opcodes_h_l652_c2_885b_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_return_output := t16_MUX_uxn_opcodes_h_l652_c2_885b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l652_c2_885b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_return_output := result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l652_c2_885b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output;

     -- Submodule level 7
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l652_c2_885b_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l681_l648_DUPLICATE_1d01 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l681_l648_DUPLICATE_1d01_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l652_c2_885b_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l681_l648_DUPLICATE_1d01_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_cc5c_uxn_opcodes_h_l681_l648_DUPLICATE_1d01_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
