-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity gth_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_6d7675a8;
architecture arch of gth_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1916_c6_ee4c]
signal BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1916_c1_522c]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1916_c2_1754]
signal n8_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1916_c2_1754]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1916_c2_1754]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1916_c2_1754]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1916_c2_1754]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1916_c2_1754]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1916_c2_1754]
signal result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1916_c2_1754]
signal t8_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1917_c3_70aa[uxn_opcodes_h_l1917_c3_70aa]
signal printf_uxn_opcodes_h_l1917_c3_70aa_uxn_opcodes_h_l1917_c3_70aa_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1921_c11_e71a]
signal BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1921_c7_5d04]
signal n8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1921_c7_5d04]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1921_c7_5d04]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1921_c7_5d04]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1921_c7_5d04]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1921_c7_5d04]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1921_c7_5d04]
signal result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1921_c7_5d04]
signal t8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1924_c11_7d06]
signal BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1924_c7_4b23]
signal n8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1924_c7_4b23]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1924_c7_4b23]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1924_c7_4b23]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1924_c7_4b23]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1924_c7_4b23]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1924_c7_4b23]
signal result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1924_c7_4b23]
signal t8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1928_c11_8e4b]
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1928_c7_eff5]
signal n8_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1928_c7_eff5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1928_c7_eff5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1928_c7_eff5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1928_c7_eff5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1928_c7_eff5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1928_c7_eff5]
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1931_c11_491f]
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1931_c7_172f]
signal n8_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1931_c7_172f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1931_c7_172f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1931_c7_172f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1931_c7_172f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1931_c7_172f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1931_c7_172f]
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1934_c30_3c8b]
signal sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1937_c21_4607]
signal BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1937_c21_7057]
signal MUX_uxn_opcodes_h_l1937_c21_7057_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1937_c21_7057_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1937_c21_7057_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1937_c21_7057_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1939_c11_9839]
signal BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1939_c7_1bd5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1939_c7_1bd5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1939_c7_1bd5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c
BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_left,
BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_right,
BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_return_output);

-- n8_MUX_uxn_opcodes_h_l1916_c2_1754
n8_MUX_uxn_opcodes_h_l1916_c2_1754 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1916_c2_1754_cond,
n8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue,
n8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse,
n8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754
result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754
result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754
result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754
result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754
result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_cond,
result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

-- t8_MUX_uxn_opcodes_h_l1916_c2_1754
t8_MUX_uxn_opcodes_h_l1916_c2_1754 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1916_c2_1754_cond,
t8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue,
t8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse,
t8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

-- printf_uxn_opcodes_h_l1917_c3_70aa_uxn_opcodes_h_l1917_c3_70aa
printf_uxn_opcodes_h_l1917_c3_70aa_uxn_opcodes_h_l1917_c3_70aa : entity work.printf_uxn_opcodes_h_l1917_c3_70aa_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1917_c3_70aa_uxn_opcodes_h_l1917_c3_70aa_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a
BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_left,
BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_right,
BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output);

-- n8_MUX_uxn_opcodes_h_l1921_c7_5d04
n8_MUX_uxn_opcodes_h_l1921_c7_5d04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond,
n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue,
n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse,
n8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04
result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_cond,
result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output);

-- t8_MUX_uxn_opcodes_h_l1921_c7_5d04
t8_MUX_uxn_opcodes_h_l1921_c7_5d04 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond,
t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue,
t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse,
t8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06
BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_left,
BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_right,
BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output);

-- n8_MUX_uxn_opcodes_h_l1924_c7_4b23
n8_MUX_uxn_opcodes_h_l1924_c7_4b23 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond,
n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue,
n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse,
n8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_cond,
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output);

-- t8_MUX_uxn_opcodes_h_l1924_c7_4b23
t8_MUX_uxn_opcodes_h_l1924_c7_4b23 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond,
t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue,
t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse,
t8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_left,
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_right,
BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output);

-- n8_MUX_uxn_opcodes_h_l1928_c7_eff5
n8_MUX_uxn_opcodes_h_l1928_c7_eff5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1928_c7_eff5_cond,
n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue,
n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse,
n8_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5
result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_left,
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_right,
BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output);

-- n8_MUX_uxn_opcodes_h_l1931_c7_172f
n8_MUX_uxn_opcodes_h_l1931_c7_172f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1931_c7_172f_cond,
n8_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue,
n8_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse,
n8_MUX_uxn_opcodes_h_l1931_c7_172f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_cond,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b
sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_ins,
sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_x,
sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_y,
sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607
BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607 : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_left,
BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_right,
BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_return_output);

-- MUX_uxn_opcodes_h_l1937_c21_7057
MUX_uxn_opcodes_h_l1937_c21_7057 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1937_c21_7057_cond,
MUX_uxn_opcodes_h_l1937_c21_7057_iftrue,
MUX_uxn_opcodes_h_l1937_c21_7057_iffalse,
MUX_uxn_opcodes_h_l1937_c21_7057_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839
BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_left,
BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_right,
BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5
result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5
result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5
result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_return_output,
 n8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
 t8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output,
 n8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output,
 t8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output,
 n8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output,
 t8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output,
 n8_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output,
 n8_MUX_uxn_opcodes_h_l1931_c7_172f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_return_output,
 sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_return_output,
 MUX_uxn_opcodes_h_l1937_c21_7057_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1918_c3_7416 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1917_c3_70aa_uxn_opcodes_h_l1917_c3_70aa_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_1234 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_be54 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_1dbb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1936_c3_2abf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1931_c7_172f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1937_c21_7057_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1937_c21_7057_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1937_c21_7057_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1937_c21_7057_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_2613_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_6ecf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_8f64_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_5e9e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1921_l1939_l1931_l1928_l1924_DUPLICATE_145a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1945_l1912_DUPLICATE_c80d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1936_c3_2abf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1936_c3_2abf;
     VAR_MUX_uxn_opcodes_h_l1937_c21_7057_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_1dbb := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_1dbb;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_1234 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1922_c3_1234;
     VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1918_c3_7416 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1918_c3_7416;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1937_c21_7057_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_be54 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1926_c3_be54;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_8f64 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_8f64_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1921_c11_e71a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1916_c6_ee4c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1928_c11_8e4b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1921_l1939_l1931_l1928_l1924_DUPLICATE_145a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1921_l1939_l1931_l1928_l1924_DUPLICATE_145a_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1939_c11_9839] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_left;
     BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output := BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1937_c21_4607] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_left;
     BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_return_output := BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1924_c11_7d06] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_left;
     BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output := BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_5e9e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_5e9e_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_2613 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_2613_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1931_c7_172f] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1931_c7_172f_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_6ecf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_6ecf_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1934_c30_3c8b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_ins;
     sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_x;
     sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_return_output := sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1931_c11_491f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1916_c6_ee4c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c11_e71a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1924_c11_7d06_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1928_c11_8e4b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1931_c11_491f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1939_c11_9839_return_output;
     VAR_MUX_uxn_opcodes_h_l1937_c21_7057_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1937_c21_4607_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_2613_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_2613_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_2613_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_2613_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_2613_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1921_l1939_l1931_l1928_l1924_DUPLICATE_145a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1921_l1939_l1931_l1928_l1924_DUPLICATE_145a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1921_l1939_l1931_l1928_l1924_DUPLICATE_145a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1921_l1939_l1931_l1928_l1924_DUPLICATE_145a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1921_l1939_l1931_l1928_l1924_DUPLICATE_145a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_6ecf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_6ecf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_6ecf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_6ecf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_6ecf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_8f64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_8f64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_8f64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_8f64_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1921_l1916_l1939_l1928_l1924_DUPLICATE_8f64_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_5e9e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_5e9e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_5e9e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_5e9e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1921_l1916_l1931_l1928_l1924_DUPLICATE_5e9e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1931_c7_172f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1934_c30_3c8b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1939_c7_1bd5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output;

     -- MUX[uxn_opcodes_h_l1937_c21_7057] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1937_c21_7057_cond <= VAR_MUX_uxn_opcodes_h_l1937_c21_7057_cond;
     MUX_uxn_opcodes_h_l1937_c21_7057_iftrue <= VAR_MUX_uxn_opcodes_h_l1937_c21_7057_iftrue;
     MUX_uxn_opcodes_h_l1937_c21_7057_iffalse <= VAR_MUX_uxn_opcodes_h_l1937_c21_7057_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1937_c21_7057_return_output := MUX_uxn_opcodes_h_l1937_c21_7057_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1916_c1_522c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1931_c7_172f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1931_c7_172f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1924_c7_4b23] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond <= VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond;
     t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue;
     t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output := t8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;

     -- n8_MUX[uxn_opcodes_h_l1931_c7_172f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1931_c7_172f_cond <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_cond;
     n8_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue;
     n8_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_return_output := n8_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1939_c7_1bd5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1939_c7_1bd5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue := VAR_MUX_uxn_opcodes_h_l1937_c21_7057_return_output;
     VAR_printf_uxn_opcodes_h_l1917_c3_70aa_uxn_opcodes_h_l1917_c3_70aa_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1916_c1_522c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1939_c7_1bd5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;
     -- printf_uxn_opcodes_h_l1917_c3_70aa[uxn_opcodes_h_l1917_c3_70aa] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1917_c3_70aa_uxn_opcodes_h_l1917_c3_70aa_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1917_c3_70aa_uxn_opcodes_h_l1917_c3_70aa_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1931_c7_172f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1928_c7_eff5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1928_c7_eff5] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1928_c7_eff5_cond <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_cond;
     n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue;
     n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output := n8_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1931_c7_172f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_return_output := result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1931_c7_172f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1931_c7_172f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;

     -- t8_MUX[uxn_opcodes_h_l1921_c7_5d04] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond <= VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond;
     t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue;
     t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output := t8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1928_c7_eff5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1931_c7_172f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;
     -- t8_MUX[uxn_opcodes_h_l1916_c2_1754] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1916_c2_1754_cond <= VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_cond;
     t8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue;
     t8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output := t8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1928_c7_eff5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;

     -- n8_MUX[uxn_opcodes_h_l1924_c7_4b23] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond <= VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_cond;
     n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue;
     n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output := n8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1924_c7_4b23] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1928_c7_eff5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1928_c7_eff5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1928_c7_eff5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1924_c7_4b23] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1928_c7_eff5_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1924_c7_4b23] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1924_c7_4b23] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1921_c7_5d04] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;

     -- n8_MUX[uxn_opcodes_h_l1921_c7_5d04] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond <= VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_cond;
     n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue;
     n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output := n8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1921_c7_5d04] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1924_c7_4b23] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1924_c7_4b23] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output := result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1924_c7_4b23_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1921_c7_5d04] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1921_c7_5d04] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1916_c2_1754] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1921_c7_5d04] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1921_c7_5d04] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output := result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;

     -- n8_MUX[uxn_opcodes_h_l1916_c2_1754] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1916_c2_1754_cond <= VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_cond;
     n8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue;
     n8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output := n8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1916_c2_1754] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c7_5d04_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1916_c2_1754] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1916_c2_1754] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1916_c2_1754] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1916_c2_1754] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_return_output := result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1945_l1912_DUPLICATE_c80d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1945_l1912_DUPLICATE_c80d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1916_c2_1754_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1916_c2_1754_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1945_l1912_DUPLICATE_c80d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l1945_l1912_DUPLICATE_c80d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
