-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity ldz_0CLK_46731a7b is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_46731a7b;
architecture arch of ldz_0CLK_46731a7b is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1518_c6_b4b2]
signal BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1518_c1_2144]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1518_c2_2832]
signal tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1518_c2_2832]
signal t8_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1518_c2_2832]
signal result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1518_c2_2832]
signal result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1518_c2_2832]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1518_c2_2832]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1518_c2_2832]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1518_c2_2832]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1518_c2_2832]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(3 downto 0);

-- printf_uxn_opcodes_h_l1519_c3_6f36[uxn_opcodes_h_l1519_c3_6f36]
signal printf_uxn_opcodes_h_l1519_c3_6f36_uxn_opcodes_h_l1519_c3_6f36_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1523_c11_9403]
signal BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1523_c7_ba8b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1526_c11_c4db]
signal BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1526_c7_553c]
signal tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1526_c7_553c]
signal t8_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1526_c7_553c]
signal result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1526_c7_553c]
signal result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1526_c7_553c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1526_c7_553c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1526_c7_553c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1526_c7_553c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1526_c7_553c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1529_c30_d90a]
signal sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1532_c11_b34c]
signal BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1532_c7_7821]
signal tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1532_c7_7821]
signal result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1532_c7_7821]
signal result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1532_c7_7821]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1532_c7_7821]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1532_c7_7821]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1532_c7_7821]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1536_c11_e28d]
signal BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1536_c7_5ee5]
signal tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1536_c7_5ee5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1536_c7_5ee5]
signal result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1536_c7_5ee5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1536_c7_5ee5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1542_c11_bed4]
signal BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1542_c7_8619]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1542_c7_8619]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_9969( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.u16_value := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2
BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_left,
BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_right,
BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1518_c2_2832
tmp8_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- t8_MUX_uxn_opcodes_h_l1518_c2_2832
t8_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
t8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
t8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
t8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832
result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832
result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832
result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832
result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832
result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832
result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

-- printf_uxn_opcodes_h_l1519_c3_6f36_uxn_opcodes_h_l1519_c3_6f36
printf_uxn_opcodes_h_l1519_c3_6f36_uxn_opcodes_h_l1519_c3_6f36 : entity work.printf_uxn_opcodes_h_l1519_c3_6f36_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1519_c3_6f36_uxn_opcodes_h_l1519_c3_6f36_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403
BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_left,
BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_right,
BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b
tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- t8_MUX_uxn_opcodes_h_l1523_c7_ba8b
t8_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b
result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b
result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db
BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_left,
BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_right,
BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1526_c7_553c
tmp8_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- t8_MUX_uxn_opcodes_h_l1526_c7_553c
t8_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
t8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
t8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
t8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a
sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_ins,
sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_x,
sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_y,
sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c
BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_left,
BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_right,
BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1532_c7_7821
tmp8_MUX_uxn_opcodes_h_l1532_c7_7821 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_cond,
tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue,
tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse,
tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond,
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond,
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d
BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_left,
BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_right,
BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5
tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond,
tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue,
tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse,
tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5
result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond,
result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4
BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_left,
BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_right,
BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_return_output,
 tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 t8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output,
 tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output,
 tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 t8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output,
 tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output,
 tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iffalse : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1520_c3_0637 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1519_c3_6f36_uxn_opcodes_h_l1519_c3_6f36_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1524_c3_77bf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1530_c22_d8e7_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1534_c22_6a32_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1539_c3_5e86 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1536_DUPLICATE_be4b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_38a2_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1518_l1523_l1526_DUPLICATE_51f4_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1542_DUPLICATE_d45e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_5ab4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1542_l1536_DUPLICATE_8a57_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1532_l1536_l1526_DUPLICATE_c956_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1547_l1514_DUPLICATE_a5ee_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1520_c3_0637 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1520_c3_0637;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_right := to_unsigned(5, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1524_c3_77bf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1524_c3_77bf;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1539_c3_5e86 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1539_c3_5e86;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse := tmp8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1523_c11_9403] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_left;
     BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output := BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1536_c11_e28d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1526_c11_c4db] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_left;
     BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output := BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1542_c11_bed4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1518_c6_b4b2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1542_l1536_DUPLICATE_8a57 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1542_l1536_DUPLICATE_8a57_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_38a2 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_38a2_return_output := result.u16_value;

     -- sp_relative_shift[uxn_opcodes_h_l1529_c30_d90a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_ins;
     sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_x;
     sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_return_output := sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1534_c22_6a32] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1534_c22_6a32_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1536_DUPLICATE_be4b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1536_DUPLICATE_be4b_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1518_l1523_l1526_DUPLICATE_51f4 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1518_l1523_l1526_DUPLICATE_51f4_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_5ab4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_5ab4_return_output := result.is_sp_shift;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1530_c22_d8e7] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1530_c22_d8e7_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1532_l1536_l1526_DUPLICATE_c956 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1532_l1536_l1526_DUPLICATE_c956_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1532_c11_b34c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1542_DUPLICATE_d45e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1542_DUPLICATE_d45e_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1518_c6_b4b2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1523_c11_9403_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1526_c11_c4db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1532_c11_b34c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1536_c11_e28d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1542_c11_bed4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1530_c22_d8e7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1534_c22_6a32_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1518_l1523_l1526_DUPLICATE_51f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1518_l1523_l1526_DUPLICATE_51f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1518_l1523_l1526_DUPLICATE_51f4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_38a2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_38a2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_38a2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1542_l1536_DUPLICATE_8a57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1542_l1536_DUPLICATE_8a57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1542_l1536_DUPLICATE_8a57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1542_l1536_DUPLICATE_8a57_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1542_l1536_DUPLICATE_8a57_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_5ab4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_5ab4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1518_l1532_l1523_DUPLICATE_5ab4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1542_DUPLICATE_d45e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1542_DUPLICATE_d45e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1542_DUPLICATE_d45e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1542_DUPLICATE_d45e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1542_DUPLICATE_d45e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1532_l1536_l1526_DUPLICATE_c956_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1532_l1536_l1526_DUPLICATE_c956_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1532_l1536_l1526_DUPLICATE_c956_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1536_DUPLICATE_be4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1536_DUPLICATE_be4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1536_DUPLICATE_be4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1536_DUPLICATE_be4b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1532_l1526_l1523_l1518_l1536_DUPLICATE_be4b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1529_c30_d90a_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1536_c7_5ee5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1542_c7_8619] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1542_c7_8619] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_return_output;

     -- t8_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     t8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     t8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := t8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1532_c7_7821] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output := result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1536_c7_5ee5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output := result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1518_c1_2144] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1536_c7_5ee5] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond;
     tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output := tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1532_c7_7821] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l1519_c3_6f36_uxn_opcodes_h_l1519_c3_6f36_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1518_c1_2144_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1542_c7_8619_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1542_c7_8619_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;
     -- printf_uxn_opcodes_h_l1519_c3_6f36[uxn_opcodes_h_l1519_c3_6f36] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1519_c3_6f36_uxn_opcodes_h_l1519_c3_6f36_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1519_c3_6f36_uxn_opcodes_h_l1519_c3_6f36_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1532_c7_7821] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1532_c7_7821] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output := result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- t8_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1536_c7_5ee5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1536_c7_5ee5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1532_c7_7821] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_cond;
     tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_return_output := tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1536_c7_5ee5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1532_c7_7821] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;

     -- t8_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     t8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     t8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := t8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1532_c7_7821] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1532_c7_7821_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1526_c7_553c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1526_c7_553c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1523_c7_ba8b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1523_c7_ba8b_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1518_c2_2832] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1547_l1514_DUPLICATE_a5ee LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1547_l1514_DUPLICATE_a5ee_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_9969(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1518_c2_2832_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1518_c2_2832_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1547_l1514_DUPLICATE_a5ee_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9969_uxn_opcodes_h_l1547_l1514_DUPLICATE_a5ee_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
