-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2640_c6_2285]
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal n8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal l8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2640_c2_16c1]
signal t8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2653_c11_2e4e]
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2653_c7_3001]
signal n8_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2653_c7_3001]
signal l8_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2653_c7_3001]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2653_c7_3001]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2653_c7_3001]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2653_c7_3001]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2653_c7_3001]
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2653_c7_3001]
signal t8_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2656_c11_e258]
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2656_c7_8783]
signal n8_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2656_c7_8783]
signal l8_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c7_8783]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c7_8783]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c7_8783]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c7_8783]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2656_c7_8783]
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2656_c7_8783]
signal t8_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2660_c11_90dc]
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2660_c7_3eaf]
signal n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2660_c7_3eaf]
signal l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2660_c7_3eaf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2660_c7_3eaf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2660_c7_3eaf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2660_c7_3eaf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2660_c7_3eaf]
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2662_c30_e290]
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2667_c11_8097]
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2667_c7_04e5]
signal l8_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2667_c7_04e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2667_c7_04e5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2667_c7_04e5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2667_c7_04e5]
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_561f]
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_4313]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_4313]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_4313]
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_04b4( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_vram_write := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_left,
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_right,
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output);

-- n8_MUX_uxn_opcodes_h_l2640_c2_16c1
n8_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
n8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- l8_MUX_uxn_opcodes_h_l2640_c2_16c1
l8_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
l8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- t8_MUX_uxn_opcodes_h_l2640_c2_16c1
t8_MUX_uxn_opcodes_h_l2640_c2_16c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond,
t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue,
t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse,
t8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_left,
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_right,
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output);

-- n8_MUX_uxn_opcodes_h_l2653_c7_3001
n8_MUX_uxn_opcodes_h_l2653_c7_3001 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2653_c7_3001_cond,
n8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue,
n8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse,
n8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output);

-- l8_MUX_uxn_opcodes_h_l2653_c7_3001
l8_MUX_uxn_opcodes_h_l2653_c7_3001 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2653_c7_3001_cond,
l8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue,
l8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse,
l8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_cond,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_return_output);

-- t8_MUX_uxn_opcodes_h_l2653_c7_3001
t8_MUX_uxn_opcodes_h_l2653_c7_3001 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2653_c7_3001_cond,
t8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue,
t8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse,
t8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_left,
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_right,
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output);

-- n8_MUX_uxn_opcodes_h_l2656_c7_8783
n8_MUX_uxn_opcodes_h_l2656_c7_8783 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2656_c7_8783_cond,
n8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue,
n8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse,
n8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output);

-- l8_MUX_uxn_opcodes_h_l2656_c7_8783
l8_MUX_uxn_opcodes_h_l2656_c7_8783 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2656_c7_8783_cond,
l8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue,
l8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse,
l8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_cond,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_return_output);

-- t8_MUX_uxn_opcodes_h_l2656_c7_8783
t8_MUX_uxn_opcodes_h_l2656_c7_8783 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2656_c7_8783_cond,
t8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue,
t8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse,
t8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_left,
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_right,
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output);

-- n8_MUX_uxn_opcodes_h_l2660_c7_3eaf
n8_MUX_uxn_opcodes_h_l2660_c7_3eaf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond,
n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue,
n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse,
n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output);

-- l8_MUX_uxn_opcodes_h_l2660_c7_3eaf
l8_MUX_uxn_opcodes_h_l2660_c7_3eaf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond,
l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue,
l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse,
l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2662_c30_e290
sp_relative_shift_uxn_opcodes_h_l2662_c30_e290 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_ins,
sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_x,
sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_y,
sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_left,
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_right,
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output);

-- l8_MUX_uxn_opcodes_h_l2667_c7_04e5
l8_MUX_uxn_opcodes_h_l2667_c7_04e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2667_c7_04e5_cond,
l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue,
l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse,
l8_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_cond,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_left,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_right,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_cond,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output,
 n8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 l8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 t8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output,
 n8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output,
 l8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_return_output,
 t8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output,
 n8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output,
 l8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_return_output,
 t8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output,
 n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output,
 l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output,
 sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output,
 l8_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_8927 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_937f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_6aa6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_d55b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_818c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_19d1 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_f462 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_1209 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_4313_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_3074_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_09ca_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2660_l2656_l2653_l2673_l2667_DUPLICATE_2a56_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_c6f3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2679_l2636_DUPLICATE_e6e3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_19d1 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_19d1;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_6aa6 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_6aa6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_8927 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_8927;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_818c := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_818c;
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_1209 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_1209;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_f462 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_f462;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_937f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_937f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_d55b := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_d55b;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse := t8;
     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_09ca LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_09ca_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2660_l2656_l2653_l2673_l2667_DUPLICATE_2a56 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2660_l2656_l2653_l2673_l2667_DUPLICATE_2a56_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2656_c11_e258] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_left;
     BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output := BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2640_c6_2285] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_left;
     BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output := BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2660_c11_90dc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_left;
     BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output := BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2653_c11_2e4e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2662_c30_e290] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_ins;
     sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_x;
     sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_return_output := sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_561f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output := result.is_vram_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2673_c7_4313] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_4313_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_3074 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_3074_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2667_c11_8097] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_left;
     BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output := BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_c6f3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_c6f3_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_2285_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_2e4e_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_e258_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_90dc_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_8097_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_561f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_09ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_09ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_09ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2660_l2656_l2653_l2673_l2667_DUPLICATE_2a56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2660_l2656_l2653_l2673_l2667_DUPLICATE_2a56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2660_l2656_l2653_l2673_l2667_DUPLICATE_2a56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2660_l2656_l2653_l2673_l2667_DUPLICATE_2a56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2660_l2656_l2653_l2673_l2667_DUPLICATE_2a56_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_c6f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_c6f3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2660_l2653_l2656_DUPLICATE_c6f3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_3074_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_3074_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_3074_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2673_l2640_l2653_l2656_DUPLICATE_3074_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_16c1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_4313_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_e290_return_output;
     -- n8_MUX[uxn_opcodes_h_l2660_c7_3eaf] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond;
     n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue;
     n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output := n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2667_c7_04e5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_4313] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- t8_MUX[uxn_opcodes_h_l2656_c7_8783] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2656_c7_8783_cond <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_cond;
     t8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue;
     t8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output := t8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- l8_MUX[uxn_opcodes_h_l2667_c7_04e5] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2667_c7_04e5_cond <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_cond;
     l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue;
     l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output := l8_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2660_c7_3eaf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_4313] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_4313] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_return_output := result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_4313_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_4313_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_4313_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2667_c7_04e5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;

     -- l8_MUX[uxn_opcodes_h_l2660_c7_3eaf] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond;
     l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue;
     l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output := l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;

     -- n8_MUX[uxn_opcodes_h_l2656_c7_8783] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2656_c7_8783_cond <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_cond;
     n8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue;
     n8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output := n8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2660_c7_3eaf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2667_c7_04e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c7_8783] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;

     -- t8_MUX[uxn_opcodes_h_l2653_c7_3001] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2653_c7_3001_cond <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_cond;
     t8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue;
     t8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output := t8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2667_c7_04e5] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output := result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_04e5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;
     -- l8_MUX[uxn_opcodes_h_l2656_c7_8783] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2656_c7_8783_cond <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_cond;
     l8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue;
     l8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output := l8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2660_c7_3eaf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;

     -- t8_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := t8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- n8_MUX[uxn_opcodes_h_l2653_c7_3001] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2653_c7_3001_cond <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_cond;
     n8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue;
     n8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output := n8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2660_c7_3eaf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output := result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c7_8783] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2653_c7_3001] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2660_c7_3eaf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_3eaf_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c7_8783] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;

     -- l8_MUX[uxn_opcodes_h_l2653_c7_3001] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2653_c7_3001_cond <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_cond;
     l8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue;
     l8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output := l8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2656_c7_8783] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_return_output := result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2653_c7_3001] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;

     -- n8_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := n8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c7_8783] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_8783_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2653_c7_3001] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2653_c7_3001] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_return_output := result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;

     -- l8_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := l8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2653_c7_3001] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_3001_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2640_c2_16c1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2679_l2636_DUPLICATE_e6e3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2679_l2636_DUPLICATE_e6e3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_04b4(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_16c1_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2679_l2636_DUPLICATE_e6e3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_04b4_uxn_opcodes_h_l2679_l2636_DUPLICATE_e6e3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
