-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 57
entity mul_0CLK_edc09f97 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_edc09f97;
architecture arch of mul_0CLK_edc09f97 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2139_c6_6df6]
signal BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2139_c2_153c]
signal n8_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2139_c2_153c]
signal t8_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2139_c2_153c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2139_c2_153c]
signal result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2139_c2_153c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2139_c2_153c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2139_c2_153c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2139_c2_153c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2144_c11_6884]
signal BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2144_c7_7989]
signal n8_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2144_c7_7989]
signal t8_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2144_c7_7989]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2144_c7_7989]
signal result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2144_c7_7989]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2144_c7_7989]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2144_c7_7989]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2144_c7_7989]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2147_c11_7d04]
signal BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2147_c7_09fa]
signal n8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2147_c7_09fa]
signal t8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2147_c7_09fa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2147_c7_09fa]
signal result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2147_c7_09fa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2147_c7_09fa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2147_c7_09fa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2147_c7_09fa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2151_c11_e079]
signal BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2151_c7_70cd]
signal n8_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2151_c7_70cd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2151_c7_70cd]
signal result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2151_c7_70cd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2151_c7_70cd]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2151_c7_70cd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2151_c7_70cd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2154_c11_66fd]
signal BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2154_c7_7a17]
signal n8_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2154_c7_7a17]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2154_c7_7a17]
signal result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2154_c7_7a17]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2154_c7_7a17]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2154_c7_7a17]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2154_c7_7a17]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2157_c32_8280]
signal BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l2157_c32_968c]
signal BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2157_c32_18c9]
signal MUX_uxn_opcodes_h_l2157_c32_18c9_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2157_c32_18c9_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2157_c32_18c9_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l2157_c32_18c9_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2159_c11_3c5c]
signal BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l2159_c7_f203]
signal result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2159_c7_f203]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2159_c7_f203]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2159_c7_f203]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2159_c7_f203]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(0 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2163_c24_310b]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2165_c11_6552]
signal BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2165_c7_313b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2165_c7_313b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.is_opc_done := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6
BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_left,
BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_right,
BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output);

-- n8_MUX_uxn_opcodes_h_l2139_c2_153c
n8_MUX_uxn_opcodes_h_l2139_c2_153c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2139_c2_153c_cond,
n8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue,
n8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse,
n8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

-- t8_MUX_uxn_opcodes_h_l2139_c2_153c
t8_MUX_uxn_opcodes_h_l2139_c2_153c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2139_c2_153c_cond,
t8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue,
t8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse,
t8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c
result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_cond,
result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c
result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c
result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c
result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884
BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_left,
BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_right,
BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output);

-- n8_MUX_uxn_opcodes_h_l2144_c7_7989
n8_MUX_uxn_opcodes_h_l2144_c7_7989 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2144_c7_7989_cond,
n8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue,
n8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse,
n8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output);

-- t8_MUX_uxn_opcodes_h_l2144_c7_7989
t8_MUX_uxn_opcodes_h_l2144_c7_7989 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2144_c7_7989_cond,
t8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue,
t8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse,
t8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989
result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_cond,
result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989
result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04
BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_left,
BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_right,
BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output);

-- n8_MUX_uxn_opcodes_h_l2147_c7_09fa
n8_MUX_uxn_opcodes_h_l2147_c7_09fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond,
n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue,
n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse,
n8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output);

-- t8_MUX_uxn_opcodes_h_l2147_c7_09fa
t8_MUX_uxn_opcodes_h_l2147_c7_09fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond,
t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue,
t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse,
t8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa
result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_cond,
result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa
result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079
BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_left,
BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_right,
BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output);

-- n8_MUX_uxn_opcodes_h_l2151_c7_70cd
n8_MUX_uxn_opcodes_h_l2151_c7_70cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2151_c7_70cd_cond,
n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue,
n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse,
n8_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd
result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_cond,
result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd
result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd
BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_left,
BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_right,
BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output);

-- n8_MUX_uxn_opcodes_h_l2154_c7_7a17
n8_MUX_uxn_opcodes_h_l2154_c7_7a17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2154_c7_7a17_cond,
n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue,
n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse,
n8_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17
result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17
result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_cond,
result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17
result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17
result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17
result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280
BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_left,
BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_right,
BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c
BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_left,
BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_right,
BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_return_output);

-- MUX_uxn_opcodes_h_l2157_c32_18c9
MUX_uxn_opcodes_h_l2157_c32_18c9 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2157_c32_18c9_cond,
MUX_uxn_opcodes_h_l2157_c32_18c9_iftrue,
MUX_uxn_opcodes_h_l2157_c32_18c9_iffalse,
MUX_uxn_opcodes_h_l2157_c32_18c9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c
BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_left,
BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_right,
BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203
result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_cond,
result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203
result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552
BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_left,
BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_right,
BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b
result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b
result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output,
 n8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
 t8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output,
 n8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output,
 t8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output,
 n8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output,
 t8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output,
 n8_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output,
 n8_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_return_output,
 BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_return_output,
 MUX_uxn_opcodes_h_l2157_c32_18c9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2141_c3_6e62 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2145_c3_289a : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2149_c3_413d : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2152_c3_9b15 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_uxn_opcodes_h_l2163_c3_41c3 : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2162_c3_383f : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2154_l2151_l2147_l2144_l2139_DUPLICATE_6358_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2159_l2151_l2147_l2144_l2139_DUPLICATE_9f1c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2154_l2159_DUPLICATE_661d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2170_l2135_DUPLICATE_849a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_right := to_unsigned(5, 3);
     VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_iffalse := resize(to_signed(-1, 2), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2162_c3_383f := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2162_c3_383f;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2152_c3_9b15 := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2152_c3_9b15;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2145_c3_289a := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2145_c3_289a;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2149_c3_413d := resize(to_unsigned(2, 2), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2149_c3_413d;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_right := to_unsigned(128, 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_right := to_unsigned(6, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2141_c3_6e62 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2141_c3_6e62;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_left := VAR_ins;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_left := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse := t8;
     -- BIN_OP_AND[uxn_opcodes_h_l2157_c32_8280] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_left;
     BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_return_output := BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_return_output;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l2163_c24_310b] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2139_c6_6df6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0_return_output := result.stack_value;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2154_l2151_l2147_l2144_l2139_DUPLICATE_6358 LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2154_l2151_l2147_l2144_l2139_DUPLICATE_6358_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2154_l2159_DUPLICATE_661d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2154_l2159_DUPLICATE_661d_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2159_c11_3c5c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2159_l2151_l2147_l2144_l2139_DUPLICATE_9f1c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2159_l2151_l2147_l2144_l2139_DUPLICATE_9f1c_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2151_c11_e079] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_left;
     BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output := BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2144_c11_6884] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_left;
     BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output := BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2154_c11_66fd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_left;
     BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output := BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2165_c11_6552] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_left;
     BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_return_output := BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2147_c11_7d04] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_left;
     BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output := BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_left := VAR_BIN_OP_AND_uxn_opcodes_h_l2157_c32_8280_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2139_c6_6df6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2144_c11_6884_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2147_c11_7d04_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2151_c11_e079_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2154_c11_66fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2159_c11_3c5c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2165_c11_6552_return_output;
     VAR_result_stack_value_uxn_opcodes_h_l2163_c3_41c3 := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l2163_c24_310b_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2154_l2151_l2147_l2144_l2139_DUPLICATE_6358_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2154_l2151_l2147_l2144_l2139_DUPLICATE_6358_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2154_l2151_l2147_l2144_l2139_DUPLICATE_6358_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2154_l2151_l2147_l2144_l2139_DUPLICATE_6358_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2154_l2151_l2147_l2144_l2139_DUPLICATE_6358_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2165_l2159_l2154_l2151_l2147_l2144_DUPLICATE_80d0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2159_l2151_l2147_l2144_l2139_DUPLICATE_9f1c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2159_l2151_l2147_l2144_l2139_DUPLICATE_9f1c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2159_l2151_l2147_l2144_l2139_DUPLICATE_9f1c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2159_l2151_l2147_l2144_l2139_DUPLICATE_9f1c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2159_l2151_l2147_l2144_l2139_DUPLICATE_9f1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2165_l2154_l2151_l2147_l2144_l2139_DUPLICATE_3b7c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2154_l2159_DUPLICATE_661d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2154_l2159_DUPLICATE_661d_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l2159_l2154_l2151_l2147_l2144_l2139_DUPLICATE_07d0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue := VAR_result_stack_value_uxn_opcodes_h_l2163_c3_41c3;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2159_c7_f203] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2159_c7_f203] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l2157_c32_968c] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_left;
     BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_return_output := BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2165_c7_313b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2147_c7_09fa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond <= VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond;
     t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue;
     t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output := t8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2165_c7_313b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2159_c7_f203] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_return_output := result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;

     -- n8_MUX[uxn_opcodes_h_l2154_c7_7a17] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2154_c7_7a17_cond <= VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_cond;
     n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue;
     n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output := n8_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l2157_c32_968c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2165_c7_313b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2165_c7_313b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;
     -- MUX[uxn_opcodes_h_l2157_c32_18c9] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2157_c32_18c9_cond <= VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_cond;
     MUX_uxn_opcodes_h_l2157_c32_18c9_iftrue <= VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_iftrue;
     MUX_uxn_opcodes_h_l2157_c32_18c9_iffalse <= VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_return_output := MUX_uxn_opcodes_h_l2157_c32_18c9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2151_c7_70cd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2151_c7_70cd_cond <= VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_cond;
     n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue;
     n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output := n8_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2154_c7_7a17] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2159_c7_f203] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;

     -- t8_MUX[uxn_opcodes_h_l2144_c7_7989] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2144_c7_7989_cond <= VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_cond;
     t8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue;
     t8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output := t8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2154_c7_7a17] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output := result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2159_c7_f203] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2154_c7_7a17] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue := VAR_MUX_uxn_opcodes_h_l2157_c32_18c9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2159_c7_f203_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;
     -- n8_MUX[uxn_opcodes_h_l2147_c7_09fa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond <= VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_cond;
     n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue;
     n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output := n8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;

     -- t8_MUX[uxn_opcodes_h_l2139_c2_153c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2139_c2_153c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_cond;
     t8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue;
     t8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output := t8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2151_c7_70cd] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2154_c7_7a17] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2154_c7_7a17] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2154_c7_7a17] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2151_c7_70cd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2151_c7_70cd] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output := result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2154_c7_7a17_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;
     -- n8_MUX[uxn_opcodes_h_l2144_c7_7989] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2144_c7_7989_cond <= VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_cond;
     n8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue;
     n8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output := n8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2151_c7_70cd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2147_c7_09fa] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output := result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2147_c7_09fa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2151_c7_70cd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2147_c7_09fa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2151_c7_70cd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2151_c7_70cd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2147_c7_09fa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;

     -- n8_MUX[uxn_opcodes_h_l2139_c2_153c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2139_c2_153c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_cond;
     n8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue;
     n8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output := n8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2144_c7_7989] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_return_output := result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2144_c7_7989] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2144_c7_7989] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2147_c7_09fa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2147_c7_09fa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2147_c7_09fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2144_c7_7989] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2144_c7_7989] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2144_c7_7989] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l2139_c2_153c] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_cond;
     result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_return_output := result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2139_c2_153c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2139_c2_153c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;

     -- Submodule level 7
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2144_c7_7989_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2139_c2_153c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2139_c2_153c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2139_c2_153c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_return_output;

     -- Submodule level 8
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2170_l2135_DUPLICATE_849a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2170_l2135_DUPLICATE_849a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2139_c2_153c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2139_c2_153c_return_output);

     -- Submodule level 9
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2170_l2135_DUPLICATE_849a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_d2e5_uxn_opcodes_h_l2170_l2135_DUPLICATE_849a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
