-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity lit2_0CLK_d6c995e8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit2_0CLK_d6c995e8;
architecture arch of lit2_0CLK_d6c995e8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l217_c6_5fd4]
signal BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l217_c2_8039]
signal tmp16_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l217_c2_8039]
signal result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l217_c2_8039]
signal result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l217_c2_8039]
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l217_c2_8039]
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l217_c2_8039]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l217_c2_8039]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l217_c2_8039]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l226_c11_bf01]
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l226_c7_da1a]
signal tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l226_c7_da1a]
signal result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l226_c7_da1a]
signal result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l226_c7_da1a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l226_c7_da1a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l226_c7_da1a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l226_c7_da1a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l226_c7_da1a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l228_c22_fbdc]
signal BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l230_c11_e670]
signal BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l230_c7_3697]
signal tmp16_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l230_c7_3697]
signal result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l230_c7_3697]
signal result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l230_c7_3697]
signal result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l230_c7_3697]
signal result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l230_c7_3697]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l230_c7_3697]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(3 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l232_c3_1214]
signal CONST_SL_8_uxn_opcodes_h_l232_c3_1214_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l232_c3_1214_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l234_c11_c898]
signal BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output : unsigned(0 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l234_c7_4d28]
signal tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(15 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l234_c7_4d28]
signal result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l234_c7_4d28]
signal result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l234_c7_4d28]
signal result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l234_c7_4d28]
signal result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l234_c7_4d28]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l234_c7_4d28]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(3 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l235_c3_3db3]
signal BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l237_c22_1117]
signal BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l242_c11_5894]
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l242_c7_4f8a]
signal result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l242_c7_4f8a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l242_c7_4f8a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l242_c7_4f8a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l242_c7_4f8a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(3 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l245_c31_1a1f]
signal CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l247_c11_32b9]
signal BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l247_c7_f255]
signal result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l247_c7_f255]
signal result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_f68f( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_pc_updated := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4
BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_left,
BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_right,
BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output);

-- tmp16_MUX_uxn_opcodes_h_l217_c2_8039
tmp16_MUX_uxn_opcodes_h_l217_c2_8039 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l217_c2_8039_cond,
tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iftrue,
tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iffalse,
tmp16_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039
result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_cond,
result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039
result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_cond,
result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039
result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039
result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039
result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01
BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_left,
BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_right,
BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output);

-- tmp16_MUX_uxn_opcodes_h_l226_c7_da1a
tmp16_MUX_uxn_opcodes_h_l226_c7_da1a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_cond,
tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue,
tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse,
tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a
result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond,
result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a
result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond,
result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a
result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc
BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_left,
BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_right,
BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670
BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_left,
BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_right,
BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output);

-- tmp16_MUX_uxn_opcodes_h_l230_c7_3697
tmp16_MUX_uxn_opcodes_h_l230_c7_3697 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l230_c7_3697_cond,
tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iftrue,
tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iffalse,
tmp16_MUX_uxn_opcodes_h_l230_c7_3697_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697
result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_cond,
result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697
result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_cond,
result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697
result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697
result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697
result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_return_output);

-- CONST_SL_8_uxn_opcodes_h_l232_c3_1214
CONST_SL_8_uxn_opcodes_h_l232_c3_1214 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l232_c3_1214_x,
CONST_SL_8_uxn_opcodes_h_l232_c3_1214_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898
BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_left,
BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_right,
BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output);

-- tmp16_MUX_uxn_opcodes_h_l234_c7_4d28
tmp16_MUX_uxn_opcodes_h_l234_c7_4d28 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_cond,
tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue,
tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse,
tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28
result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond,
result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28
result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond,
result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28
result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28
result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28
result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3
BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_left,
BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_right,
BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117
BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117 : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_left,
BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_right,
BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894
BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_left,
BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_right,
BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a
result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_cond,
result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a
result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output);

-- CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f
CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_x,
CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9
BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_left,
BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_right,
BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255
result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255
result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output,
 tmp16_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output,
 tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output,
 tmp16_MUX_uxn_opcodes_h_l230_c7_3697_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_return_output,
 CONST_SL_8_uxn_opcodes_h_l232_c3_1214_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output,
 tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_return_output,
 BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output,
 CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l222_c3_4616 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l228_c3_e44f : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l227_c3_c74b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l226_c7_da1a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l232_c3_1214_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l232_c3_1214_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l237_c3_a8e8 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_8b11 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_return_output : unsigned(16 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_a0d0_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l244_c3_7b3e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l245_c21_a208_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_dca7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l217_l247_l242_l230_l226_DUPLICATE_01b0_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_fee2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_6846_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l247_l242_l234_l230_l226_DUPLICATE_10d0_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l235_l231_DUPLICATE_178e_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l230_l234_DUPLICATE_36d2_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f68f_uxn_opcodes_h_l212_l252_DUPLICATE_4aef_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_8b11 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_8b11;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l244_c3_7b3e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l244_c3_7b3e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l227_c3_c74b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l227_c3_c74b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l222_c3_4616 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l222_c3_4616;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_right := to_unsigned(2, 2);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_left := tmp16;
     VAR_CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse := tmp16;
     -- BIN_OP_EQ[uxn_opcodes_h_l234_c11_c898] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_left;
     BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output := BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l235_l231_DUPLICATE_178e LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l235_l231_DUPLICATE_178e_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_ram_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l217_l247_l242_l230_l226_DUPLICATE_01b0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l217_l247_l242_l230_l226_DUPLICATE_01b0_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_fee2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_fee2_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l247_c11_32b9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_left;
     BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_return_output := BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l228_c22_fbdc] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_left;
     BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_return_output := BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l237_c22_1117] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_left;
     BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_return_output := BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l242_c11_5894] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_left;
     BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output := BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l226_c7_da1a_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_dca7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_dca7_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l230_c11_e670] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_left;
     BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output := BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l226_c11_bf01] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_left;
     BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output := BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;

     -- CONST_SR_8[uxn_opcodes_h_l245_c31_1a1f] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_x <= VAR_CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_return_output := CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l230_l234_DUPLICATE_36d2 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l230_l234_DUPLICATE_36d2_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l247_l242_l234_l230_l226_DUPLICATE_10d0 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l247_l242_l234_l230_l226_DUPLICATE_10d0_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l217_c6_5fd4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_left;
     BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output := BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_6846 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_6846_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c6_5fd4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_bf01_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l230_c11_e670_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l234_c11_c898_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_5894_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l247_c11_32b9_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l228_c3_e44f := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l228_c22_fbdc_return_output, 16);
     VAR_result_u16_value_uxn_opcodes_h_l237_c3_a8e8 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l237_c22_1117_return_output, 16);
     VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l235_l231_DUPLICATE_178e_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l232_c3_1214_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l235_l231_DUPLICATE_178e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l230_l234_DUPLICATE_36d2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l230_l234_DUPLICATE_36d2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l247_l242_l234_l230_l226_DUPLICATE_10d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l247_l242_l234_l230_l226_DUPLICATE_10d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l247_l242_l234_l230_l226_DUPLICATE_10d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l247_l242_l234_l230_l226_DUPLICATE_10d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l247_l242_l234_l230_l226_DUPLICATE_10d0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_fee2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_fee2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_fee2_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_fee2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l217_l247_l242_l230_l226_DUPLICATE_01b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l217_l247_l242_l230_l226_DUPLICATE_01b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l217_l247_l242_l230_l226_DUPLICATE_01b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l217_l247_l242_l230_l226_DUPLICATE_01b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l217_l247_l242_l230_l226_DUPLICATE_01b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_6846_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_6846_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_6846_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_6846_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_dca7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_dca7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_dca7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l242_l230_l217_l226_DUPLICATE_dca7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l226_c7_da1a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue := VAR_result_u16_value_uxn_opcodes_h_l228_c3_e44f;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue := VAR_result_u16_value_uxn_opcodes_h_l237_c3_a8e8;
     -- BIN_OP_OR[uxn_opcodes_h_l235_c3_3db3] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_left;
     BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_return_output := BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l234_c7_4d28] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond;
     result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output := result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l247_c7_f255] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l245_c21_a208] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l245_c21_a208_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l245_c31_1a1f_return_output);

     -- result_is_opc_done_MUX[uxn_opcodes_h_l247_c7_f255] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l232_c3_1214] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l232_c3_1214_x <= VAR_CONST_SL_8_uxn_opcodes_h_l232_c3_1214_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l232_c3_1214_return_output := CONST_SL_8_uxn_opcodes_h_l232_c3_1214_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l242_c7_4f8a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l242_c7_4f8a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;

     -- Submodule level 2
     VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l245_c21_a208_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l232_c3_1214_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l247_c7_f255_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l247_c7_f255_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l230_c7_3697] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_cond;
     result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output := result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l234_c7_4d28] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l242_c7_4f8a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l240_c21_a0d0] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_a0d0_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l235_c3_3db3_return_output);

     -- result_is_stack_write_MUX[uxn_opcodes_h_l242_c7_4f8a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l234_c7_4d28] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l217_c2_8039] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l234_c7_4d28] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_cond;
     tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue;
     tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_return_output := tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l242_c7_4f8a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output := result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_a0d0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l242_c7_4f8a_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l230_c7_3697] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l234_c7_4d28] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l230_c7_3697] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output := result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l234_c7_4d28] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l230_c7_3697] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l230_c7_3697_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_cond;
     tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iftrue;
     tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_return_output := tmp16_MUX_uxn_opcodes_h_l230_c7_3697_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l234_c7_4d28] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_cond;
     result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output := result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l230_c7_3697_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l230_c7_3697_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l234_c7_4d28_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l230_c7_3697_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l217_c2_8039] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_cond;
     result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output := result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l230_c7_3697] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_cond;
     tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue;
     tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_return_output := tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l230_c7_3697] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_cond;
     result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output := result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l230_c7_3697] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l230_c7_3697_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l230_c7_3697_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l230_c7_3697_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l217_c2_8039] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l217_c2_8039] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l217_c2_8039_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_cond;
     tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iftrue;
     tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_return_output := tmp16_MUX_uxn_opcodes_h_l217_c2_8039_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l217_c2_8039] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l226_c7_da1a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output := result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l226_c7_da1a_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l217_c2_8039_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l217_c2_8039] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l217_c2_8039] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l217_c2_8039] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_cond;
     result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output := result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_f68f_uxn_opcodes_h_l212_l252_DUPLICATE_4aef LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f68f_uxn_opcodes_h_l212_l252_DUPLICATE_4aef_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_f68f(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l217_c2_8039_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c2_8039_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f68f_uxn_opcodes_h_l212_l252_DUPLICATE_4aef_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_f68f_uxn_opcodes_h_l212_l252_DUPLICATE_4aef_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
