-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 42
entity opc_sft_phased_0CLK_6539e591 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_sft_phased_0CLK_6539e591;
architecture arch of opc_sft_phased_0CLK_6539e591 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l1224_c6_df75]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1224_c1_b26f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1227_c7_f99c]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1224_c2_9c40]
signal t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1224_c2_9c40]
signal n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1224_c2_9c40]
signal result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l1225_c12_0cda]
signal set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1227_c11_21f7]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1227_c1_9513]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1230_c7_680e]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1227_c7_f99c]
signal t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1227_c7_f99c]
signal n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1227_c7_f99c]
signal result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l1228_c8_9236]
signal t_register_uxn_opcodes_phased_h_l1228_c8_9236_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l1228_c8_9236_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1230_c11_a067]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1230_c1_435f]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1233_c7_4197]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1230_c7_680e]
signal t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1230_c7_680e]
signal n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1230_c7_680e]
signal result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1231_c8_e4cf]
signal n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1233_c11_9829]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1233_c1_cca6]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1236_c7_d4e9]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1233_c7_4197]
signal n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1233_c7_4197]
signal result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1234_c8_91e5]
signal n_register_uxn_opcodes_phased_h_l1234_c8_91e5_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1234_c8_91e5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1236_c11_28e1]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1236_c1_d838]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1239_c7_6af0]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1236_c7_d4e9]
signal result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l1237_c3_654e]
signal set_uxn_opcodes_phased_h_l1237_c3_654e_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1237_c3_654e_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1237_c3_654e_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1237_c3_654e_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1237_c3_654e_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1237_c3_654e_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1237_c3_654e_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1239_c11_fe70]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1239_c1_6c27]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1239_c7_6af0]
signal result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_phased_h_l1240_c41_e736]
signal BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_right : unsigned(3 downto 0);
signal BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_phased_h_l1240_c34_bd16]
signal BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_phased_h_l1240_c57_cc1c]
signal CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_phased_h_l1240_c34_5789]
signal BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_return_output : unsigned(7 downto 0);

-- put_stack[uxn_opcodes_phased_h_l1240_c3_848a]
signal put_stack_uxn_opcodes_phased_h_l1240_c3_848a_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1240_c3_848a_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1240_c3_848a_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1240_c3_848a_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1240_c3_848a_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1242_c11_a584]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1242_c7_87b2]
signal result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75
BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40
t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond,
t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40
n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond,
n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40
result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond,
result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue,
result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse,
result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda
set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_sp,
set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_k,
set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_mul,
set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_add,
set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7
BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c
t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond,
t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c
n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond,
n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c
result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond,
result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue,
result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse,
result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output);

-- t_register_uxn_opcodes_phased_h_l1228_c8_9236
t_register_uxn_opcodes_phased_h_l1228_c8_9236 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l1228_c8_9236_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_index,
t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_ptr,
t_register_uxn_opcodes_phased_h_l1228_c8_9236_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067
BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e
t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond,
t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e
n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond,
n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1230_c7_680e
result_MUX_uxn_opcodes_phased_h_l1230_c7_680e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond,
result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue,
result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse,
result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output);

-- n_register_uxn_opcodes_phased_h_l1231_c8_e4cf
n_register_uxn_opcodes_phased_h_l1231_c8_e4cf : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_index,
n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_ptr,
n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829
BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197
n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond,
n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1233_c7_4197
result_MUX_uxn_opcodes_phased_h_l1233_c7_4197 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond,
result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue,
result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse,
result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output);

-- n_register_uxn_opcodes_phased_h_l1234_c8_91e5
n_register_uxn_opcodes_phased_h_l1234_c8_91e5 : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1234_c8_91e5_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_index,
n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_ptr,
n_register_uxn_opcodes_phased_h_l1234_c8_91e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1
BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9
result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond,
result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue,
result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse,
result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output);

-- set_uxn_opcodes_phased_h_l1237_c3_654e
set_uxn_opcodes_phased_h_l1237_c3_654e : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l1237_c3_654e_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l1237_c3_654e_sp,
set_uxn_opcodes_phased_h_l1237_c3_654e_stack_index,
set_uxn_opcodes_phased_h_l1237_c3_654e_ins,
set_uxn_opcodes_phased_h_l1237_c3_654e_k,
set_uxn_opcodes_phased_h_l1237_c3_654e_mul,
set_uxn_opcodes_phased_h_l1237_c3_654e_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70
BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0
result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond,
result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue,
result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse,
result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output);

-- BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736
BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736 : entity work.BIN_OP_AND_uint8_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_left,
BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_right,
BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_return_output);

-- BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16
BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16 : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_left,
BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_right,
BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_return_output);

-- CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c
CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_x,
CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_return_output);

-- BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789
BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789 : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_left,
BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_right,
BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_return_output);

-- put_stack_uxn_opcodes_phased_h_l1240_c3_848a
put_stack_uxn_opcodes_phased_h_l1240_c3_848a : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l1240_c3_848a_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l1240_c3_848a_sp,
put_stack_uxn_opcodes_phased_h_l1240_c3_848a_stack_index,
put_stack_uxn_opcodes_phased_h_l1240_c3_848a_offset,
put_stack_uxn_opcodes_phased_h_l1240_c3_848a_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584
BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2
result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_cond,
result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iftrue,
result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iffalse,
result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output,
 result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output,
 set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output,
 result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output,
 t_register_uxn_opcodes_phased_h_l1228_c8_9236_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output,
 result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output,
 n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output,
 result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output,
 n_register_uxn_opcodes_phased_h_l1234_c8_91e5_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output,
 result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_return_output,
 result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output,
 BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_return_output,
 BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_return_output,
 CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_return_output,
 BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_return_output,
 result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_value : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_return_output : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_right := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iffalse := to_unsigned(0, 1);
     VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iftrue := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_add := resize(to_signed(-1, 2), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_right := to_unsigned(2, 2);
     VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_right := to_unsigned(15, 4);
     VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_offset := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_add := resize(to_signed(-1, 2), 8);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iffalse := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_mul := resize(to_unsigned(2, 2), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_k := VAR_k;
     VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_left := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_index := VAR_stack_index;
     VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_x := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1233_c11_9829] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1230_c11_a067] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1242_c11_a584] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1236_c11_28e1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output;

     -- BIN_OP_AND[uxn_opcodes_phased_h_l1240_c41_e736] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_left <= VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_left;
     BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_right <= VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_return_output := BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1227_c11_21f7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1224_c6_df75] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1239_c11_fe70] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_return_output;

     -- CONST_SR_4[uxn_opcodes_phased_h_l1240_c57_cc1c] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_x <= VAR_CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_return_output := CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_return_output;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_right := VAR_BIN_OP_AND_uxn_opcodes_phased_h_l1240_c41_e736_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1224_c6_df75_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1227_c11_21f7_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1230_c11_a067_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1233_c11_9829_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1236_c11_28e1_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1239_c11_fe70_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1242_c11_a584_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_right := VAR_CONST_SR_4_uxn_opcodes_phased_h_l1240_c57_cc1c_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1224_c1_b26f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1242_c7_87b2] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_cond;
     result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_return_output := result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_return_output;

     -- BIN_OP_SR[uxn_opcodes_phased_h_l1240_c34_bd16] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_left <= VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_left;
     BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_right <= VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_return_output := BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1227_c7_f99c] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_left := VAR_BIN_OP_SR_uxn_opcodes_phased_h_l1240_c34_bd16_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1224_c1_b26f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1242_c7_87b2_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l1239_c7_6af0] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond;
     result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output := result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1227_c1_9513] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_return_output;

     -- BIN_OP_SL[uxn_opcodes_phased_h_l1240_c34_5789] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_left <= VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_left;
     BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_right <= VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_return_output := BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1230_c7_680e] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l1225_c12_0cda] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_sp;
     set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_k;
     set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_mul;
     set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_return_output := set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_return_output;

     -- Submodule level 3
     VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_value := VAR_BIN_OP_SL_uxn_opcodes_phased_h_l1240_c34_5789_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1227_c1_9513_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l1225_c12_0cda_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1233_c7_4197] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1236_c7_d4e9] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond;
     result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output := result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output;

     -- t_register[uxn_opcodes_phased_h_l1228_c8_9236] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l1228_c8_9236_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_index;
     t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_return_output := t_register_uxn_opcodes_phased_h_l1228_c8_9236_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1230_c1_435f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1230_c1_435f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue := VAR_t_register_uxn_opcodes_phased_h_l1228_c8_9236_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1233_c1_cca6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1236_c7_d4e9] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output;

     -- n_register[uxn_opcodes_phased_h_l1231_c8_e4cf] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_index;
     n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_return_output := n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1233_c7_4197] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond;
     result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output := result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c7_d4e9_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1233_c1_cca6_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1231_c8_e4cf_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1239_c7_6af0] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1230_c7_680e] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond;
     result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output := result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1236_c1_d838] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_return_output;

     -- n_register[uxn_opcodes_phased_h_l1234_c8_91e5] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1234_c8_91e5_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_index;
     n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_return_output := n_register_uxn_opcodes_phased_h_l1234_c8_91e5_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1230_c7_680e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond;
     t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output := t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c7_6af0_return_output;
     VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1236_c1_d838_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1234_c8_91e5_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1239_c1_6c27] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_return_output;

     -- set[uxn_opcodes_phased_h_l1237_c3_654e] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l1237_c3_654e_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l1237_c3_654e_sp <= VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_sp;
     set_uxn_opcodes_phased_h_l1237_c3_654e_stack_index <= VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_stack_index;
     set_uxn_opcodes_phased_h_l1237_c3_654e_ins <= VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_ins;
     set_uxn_opcodes_phased_h_l1237_c3_654e_k <= VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_k;
     set_uxn_opcodes_phased_h_l1237_c3_654e_mul <= VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_mul;
     set_uxn_opcodes_phased_h_l1237_c3_654e_add <= VAR_set_uxn_opcodes_phased_h_l1237_c3_654e_add;
     -- Outputs

     -- n8_MUX[uxn_opcodes_phased_h_l1233_c7_4197] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_cond;
     n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output := n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1227_c7_f99c] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond;
     result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output := result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1227_c7_f99c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond;
     t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output := t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;

     -- Submodule level 7
     VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1239_c1_6c27_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1233_c7_4197_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1230_c7_680e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_cond;
     n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output := n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;

     -- put_stack[uxn_opcodes_phased_h_l1240_c3_848a] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l1240_c3_848a_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l1240_c3_848a_sp <= VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_sp;
     put_stack_uxn_opcodes_phased_h_l1240_c3_848a_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_stack_index;
     put_stack_uxn_opcodes_phased_h_l1240_c3_848a_offset <= VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_offset;
     put_stack_uxn_opcodes_phased_h_l1240_c3_848a_value <= VAR_put_stack_uxn_opcodes_phased_h_l1240_c3_848a_value;
     -- Outputs

     -- result_MUX[uxn_opcodes_phased_h_l1224_c2_9c40] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond;
     result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output := result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1224_c2_9c40] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond;
     t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output := t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output;

     -- Submodule level 8
     VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1230_c7_680e_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1227_c7_f99c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_cond;
     n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output := n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1227_c7_f99c_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1224_c2_9c40] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_cond;
     n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output := n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l1224_c2_9c40_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
