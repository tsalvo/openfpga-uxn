-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity ovr2_0CLK_57104a4d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end ovr2_0CLK_57104a4d;
architecture arch of ovr2_0CLK_57104a4d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l336_c6_9675]
signal BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l336_c2_895b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l336_c2_895b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l336_c2_895b]
signal result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l336_c2_895b]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l336_c2_895b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l336_c2_895b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l336_c2_895b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l336_c2_895b]
signal n16_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l336_c2_895b]
signal t16_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l344_c11_8da5]
signal BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l344_c7_01c3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l344_c7_01c3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l344_c7_01c3]
signal result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l344_c7_01c3]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l344_c7_01c3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l344_c7_01c3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l344_c7_01c3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l344_c7_01c3]
signal n16_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l344_c7_01c3]
signal t16_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l347_c11_c676]
signal BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l347_c7_6944]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l347_c7_6944]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l347_c7_6944]
signal result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l347_c7_6944]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l347_c7_6944]
signal result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l347_c7_6944]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l347_c7_6944]
signal result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l347_c7_6944]
signal n16_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l347_c7_6944]
signal t16_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l350_c30_1bc1]
signal sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l355_c11_1b49]
signal BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l355_c7_a4d7]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l355_c7_a4d7]
signal result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l355_c7_a4d7]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l355_c7_a4d7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l355_c7_a4d7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l355_c7_a4d7]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l355_c7_a4d7]
signal n16_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l361_c11_22cf]
signal BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l361_c7_16ee]
signal result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(15 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l361_c7_16ee]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l361_c7_16ee]
signal result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l361_c7_16ee]
signal result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l361_c7_16ee]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l365_c11_58c5]
signal BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l365_c7_bba8]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l365_c7_bba8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l365_c7_bba8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8152( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_stack_operation_16bit := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675
BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_left,
BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_right,
BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b
result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b
result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_cond,
result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b
result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b
result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b
result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- n16_MUX_uxn_opcodes_h_l336_c2_895b
n16_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l336_c2_895b_cond,
n16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
n16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
n16_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- t16_MUX_uxn_opcodes_h_l336_c2_895b
t16_MUX_uxn_opcodes_h_l336_c2_895b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l336_c2_895b_cond,
t16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue,
t16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse,
t16_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5
BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_left,
BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_right,
BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3
result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3
result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3
result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3
result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3
result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- n16_MUX_uxn_opcodes_h_l344_c7_01c3
n16_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
n16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
n16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
n16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- t16_MUX_uxn_opcodes_h_l344_c7_01c3
t16_MUX_uxn_opcodes_h_l344_c7_01c3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l344_c7_01c3_cond,
t16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue,
t16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse,
t16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676
BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_left,
BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_right,
BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944
result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944
result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_cond,
result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944
result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944
result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944
result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- n16_MUX_uxn_opcodes_h_l347_c7_6944
n16_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l347_c7_6944_cond,
n16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
n16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
n16_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- t16_MUX_uxn_opcodes_h_l347_c7_6944
t16_MUX_uxn_opcodes_h_l347_c7_6944 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l347_c7_6944_cond,
t16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue,
t16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse,
t16_MUX_uxn_opcodes_h_l347_c7_6944_return_output);

-- sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1
sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_ins,
sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_x,
sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_y,
sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49
BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_left,
BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_right,
BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7
result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7
result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_cond,
result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7
result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7
result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output);

-- n16_MUX_uxn_opcodes_h_l355_c7_a4d7
n16_MUX_uxn_opcodes_h_l355_c7_a4d7 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l355_c7_a4d7_cond,
n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue,
n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse,
n16_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf
BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_left,
BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_right,
BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee
result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_cond,
result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee
result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee
result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5
BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_left,
BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_right,
BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8
result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8
result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 n16_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 t16_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 n16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 t16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 n16_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 t16_MUX_uxn_opcodes_h_l347_c7_6944_return_output,
 sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output,
 n16_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l341_c3_c9e9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l345_c3_1b7d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l352_c3_642b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l358_c3_5c21 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l362_c3_a6bc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l361_c7_16ee_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l336_l355_l344_DUPLICATE_a10d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l336_l344_l361_DUPLICATE_51e0_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l336_l344_l347_DUPLICATE_137b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l355_l344_l336_l365_l361_DUPLICATE_c2cc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_8eab_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_eb0a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l371_l332_DUPLICATE_a2f5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_right := to_unsigned(5, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l352_c3_642b := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l352_c3_642b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l362_c3_a6bc := resize(to_unsigned(6, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l362_c3_a6bc;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l341_c3_c9e9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l341_c3_c9e9;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l345_c3_1b7d := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l345_c3_1b7d;
     VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_y := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l358_c3_5c21 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l358_c3_5c21;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse := n16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_left := VAR_phase;
     VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := t16;
     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l336_l344_l361_DUPLICATE_51e0 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l336_l344_l361_DUPLICATE_51e0_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_8eab LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_8eab_return_output := result.is_stack_operation_16bit;

     -- BIN_OP_EQ[uxn_opcodes_h_l344_c11_8da5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_left;
     BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output := BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l336_l344_l347_DUPLICATE_137b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l336_l344_l347_DUPLICATE_137b_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l361_c11_22cf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_left;
     BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output := BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_eb0a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_eb0a_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l350_c30_1bc1] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_ins;
     sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_x <= VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_x;
     sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_y <= VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_return_output := sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l336_c6_9675] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_left;
     BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output := BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l361_c7_16ee] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l361_c7_16ee_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l355_c11_1b49] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_left;
     BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output := BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l365_c11_58c5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_left;
     BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output := BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l347_c11_c676] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_left;
     BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output := BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l355_l344_l336_l365_l361_DUPLICATE_c2cc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l355_l344_l336_l365_l361_DUPLICATE_c2cc_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l336_l355_l344_DUPLICATE_a10d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l336_l355_l344_DUPLICATE_a10d_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l336_c6_9675_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l344_c11_8da5_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l347_c11_c676_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l355_c11_1b49_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l361_c11_22cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l365_c11_58c5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l336_l344_l347_DUPLICATE_137b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l336_l344_l347_DUPLICATE_137b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l336_l344_l347_DUPLICATE_137b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l336_l344_l361_DUPLICATE_51e0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l336_l344_l361_DUPLICATE_51e0_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l336_l344_l361_DUPLICATE_51e0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_eb0a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_eb0a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_eb0a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_eb0a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_eb0a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l336_l355_l344_DUPLICATE_a10d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l336_l355_l344_DUPLICATE_a10d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l336_l355_l344_DUPLICATE_a10d_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_8eab_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_8eab_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_8eab_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_8eab_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l355_l347_l344_l365_l361_DUPLICATE_8eab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l355_l344_l336_l365_l361_DUPLICATE_c2cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l355_l344_l336_l365_l361_DUPLICATE_c2cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l355_l344_l336_l365_l361_DUPLICATE_c2cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l355_l344_l336_l365_l361_DUPLICATE_c2cc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l355_l344_l336_l365_l361_DUPLICATE_c2cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l361_c7_16ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l350_c30_1bc1_return_output;
     -- n16_MUX[uxn_opcodes_h_l355_c7_a4d7] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l355_c7_a4d7_cond <= VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_cond;
     n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue;
     n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output := n16_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l365_c7_bba8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l365_c7_bba8] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l365_c7_bba8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l355_c7_a4d7] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l361_c7_16ee] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;

     -- t16_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     t16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     t16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_return_output := t16_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l361_c7_16ee] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_cond;
     result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_return_output := result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;

     -- Submodule level 2
     VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := VAR_n16_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l365_c7_bba8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l365_c7_bba8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l365_c7_bba8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_t16_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l361_c7_16ee] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l355_c7_a4d7] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l361_c7_16ee] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l361_c7_16ee] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- t16_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     t16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     t16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := t16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- n16_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     n16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     n16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_return_output := n16_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l355_c7_a4d7] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_cond;
     result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output := result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_n16_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l361_c7_16ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_t16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l355_c7_a4d7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l355_c7_a4d7] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_return_output := result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l355_c7_a4d7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- t16_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     t16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     t16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_return_output := t16_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- n16_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     n16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     n16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := n16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_n16_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l355_c7_a4d7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l336_c2_895b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- n16_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     n16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     n16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_return_output := n16_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l347_c7_6944] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l336_c2_895b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l347_c7_6944_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_return_output := result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l344_c7_01c3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l344_c7_01c3_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l336_c2_895b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l371_l332_DUPLICATE_a2f5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l371_l332_DUPLICATE_a2f5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8152(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l336_c2_895b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l336_c2_895b_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l371_l332_DUPLICATE_a2f5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8152_uxn_opcodes_h_l371_l332_DUPLICATE_a2f5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
