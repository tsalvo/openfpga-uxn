-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity sub_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_bacf6a1d;
architecture arch of sub_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2335_c6_a3a3]
signal BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2335_c1_6def]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2335_c2_443f]
signal n8_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2335_c2_443f]
signal t8_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2335_c2_443f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2335_c2_443f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2335_c2_443f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2335_c2_443f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2335_c2_443f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2335_c2_443f]
signal result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2336_c3_989a[uxn_opcodes_h_l2336_c3_989a]
signal printf_uxn_opcodes_h_l2336_c3_989a_uxn_opcodes_h_l2336_c3_989a_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2340_c11_abc4]
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2340_c7_ac3b]
signal n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2340_c7_ac3b]
signal t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2340_c7_ac3b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2340_c7_ac3b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2340_c7_ac3b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2340_c7_ac3b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2340_c7_ac3b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2340_c7_ac3b]
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2343_c11_189a]
signal BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2343_c7_3c80]
signal n8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2343_c7_3c80]
signal t8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2343_c7_3c80]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2343_c7_3c80]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2343_c7_3c80]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2343_c7_3c80]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2343_c7_3c80]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2343_c7_3c80]
signal result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2346_c11_e53c]
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2346_c7_4216]
signal n8_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2346_c7_4216]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2346_c7_4216]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2346_c7_4216]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2346_c7_4216]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2346_c7_4216]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2346_c7_4216]
signal result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2349_c30_611e]
signal sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2352_c21_8345]
signal BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2354_c11_16d1]
signal BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2354_c7_2ee8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2354_c7_2ee8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2354_c7_2ee8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3
BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_left,
BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_right,
BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_return_output);

-- n8_MUX_uxn_opcodes_h_l2335_c2_443f
n8_MUX_uxn_opcodes_h_l2335_c2_443f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2335_c2_443f_cond,
n8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue,
n8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse,
n8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

-- t8_MUX_uxn_opcodes_h_l2335_c2_443f
t8_MUX_uxn_opcodes_h_l2335_c2_443f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2335_c2_443f_cond,
t8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue,
t8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse,
t8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

-- printf_uxn_opcodes_h_l2336_c3_989a_uxn_opcodes_h_l2336_c3_989a
printf_uxn_opcodes_h_l2336_c3_989a_uxn_opcodes_h_l2336_c3_989a : entity work.printf_uxn_opcodes_h_l2336_c3_989a_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2336_c3_989a_uxn_opcodes_h_l2336_c3_989a_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_left,
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_right,
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output);

-- n8_MUX_uxn_opcodes_h_l2340_c7_ac3b
n8_MUX_uxn_opcodes_h_l2340_c7_ac3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond,
n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue,
n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse,
n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output);

-- t8_MUX_uxn_opcodes_h_l2340_c7_ac3b
t8_MUX_uxn_opcodes_h_l2340_c7_ac3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond,
t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue,
t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse,
t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a
BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_left,
BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_right,
BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output);

-- n8_MUX_uxn_opcodes_h_l2343_c7_3c80
n8_MUX_uxn_opcodes_h_l2343_c7_3c80 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond,
n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue,
n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse,
n8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output);

-- t8_MUX_uxn_opcodes_h_l2343_c7_3c80
t8_MUX_uxn_opcodes_h_l2343_c7_3c80 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond,
t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue,
t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse,
t8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_cond,
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_left,
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_right,
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output);

-- n8_MUX_uxn_opcodes_h_l2346_c7_4216
n8_MUX_uxn_opcodes_h_l2346_c7_4216 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2346_c7_4216_cond,
n8_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue,
n8_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse,
n8_MUX_uxn_opcodes_h_l2346_c7_4216_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_cond,
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2349_c30_611e
sp_relative_shift_uxn_opcodes_h_l2349_c30_611e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_ins,
sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_x,
sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_y,
sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345
BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_left,
BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_right,
BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1
BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_left,
BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_right,
BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_return_output,
 n8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
 t8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output,
 n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output,
 t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output,
 n8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output,
 t8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output,
 n8_MUX_uxn_opcodes_h_l2346_c7_4216_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_return_output,
 sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2337_c3_95f7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2336_c3_989a_uxn_opcodes_h_l2336_c3_989a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2341_c3_192f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2351_c3_1f8b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_76ba_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_71de_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_4b22_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_7493_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2346_DUPLICATE_8645_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2343_l2346_DUPLICATE_bec9_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l2360_l2331_DUPLICATE_9b98_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2351_c3_1f8b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2351_c3_1f8b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2341_c3_192f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2341_c3_192f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2337_c3_95f7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2337_c3_95f7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2340_c11_abc4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_71de LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_71de_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l2349_c30_611e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_ins;
     sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_x;
     sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_return_output := sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2352_c21_8345] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2346_c11_e53c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2346_DUPLICATE_8645 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2346_DUPLICATE_8645_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2343_c11_189a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_4b22 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_4b22_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_76ba LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_76ba_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2343_l2346_DUPLICATE_bec9 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2343_l2346_DUPLICATE_bec9_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2335_c6_a3a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_7493 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_7493_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2354_c11_16d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_a3a3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_abc4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_189a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_e53c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_16d1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_8345_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_4b22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_4b22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_4b22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_4b22_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2346_DUPLICATE_8645_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2346_DUPLICATE_8645_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2346_DUPLICATE_8645_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2346_DUPLICATE_8645_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_71de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_71de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_71de_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_71de_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_76ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_76ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_76ba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2340_l2354_l2343_l2335_DUPLICATE_76ba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2343_l2346_DUPLICATE_bec9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2343_l2346_DUPLICATE_bec9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_7493_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_7493_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_7493_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2340_l2343_l2335_l2346_DUPLICATE_7493_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_611e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2354_c7_2ee8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2335_c1_6def] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2354_c7_2ee8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2346_c7_4216] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;

     -- n8_MUX[uxn_opcodes_h_l2346_c7_4216] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2346_c7_4216_cond <= VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_cond;
     n8_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue;
     n8_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_return_output := n8_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2346_c7_4216] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2346_c7_4216] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_return_output := result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;

     -- t8_MUX[uxn_opcodes_h_l2343_c7_3c80] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond <= VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond;
     t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue;
     t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output := t8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2354_c7_2ee8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2336_c3_989a_uxn_opcodes_h_l2336_c3_989a_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_6def_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_2ee8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;
     -- t8_MUX[uxn_opcodes_h_l2340_c7_ac3b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond <= VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond;
     t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue;
     t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output := t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2343_c7_3c80] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output := result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2346_c7_4216] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2346_c7_4216] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2346_c7_4216] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;

     -- n8_MUX[uxn_opcodes_h_l2343_c7_3c80] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond <= VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_cond;
     n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue;
     n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output := n8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2343_c7_3c80] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;

     -- printf_uxn_opcodes_h_l2336_c3_989a[uxn_opcodes_h_l2336_c3_989a] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2336_c3_989a_uxn_opcodes_h_l2336_c3_989a_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2336_c3_989a_uxn_opcodes_h_l2336_c3_989a_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2343_c7_3c80] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_4216_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;
     -- n8_MUX[uxn_opcodes_h_l2340_c7_ac3b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond;
     n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue;
     n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output := n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2343_c7_3c80] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2340_c7_ac3b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2343_c7_3c80] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2340_c7_ac3b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2340_c7_ac3b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2343_c7_3c80] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;

     -- t8_MUX[uxn_opcodes_h_l2335_c2_443f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2335_c2_443f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_cond;
     t8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue;
     t8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output := t8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3c80_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;
     -- n8_MUX[uxn_opcodes_h_l2335_c2_443f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2335_c2_443f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_cond;
     n8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue;
     n8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output := n8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2335_c2_443f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2340_c7_ac3b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2340_c7_ac3b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2335_c2_443f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2340_c7_ac3b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2335_c2_443f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_ac3b_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2335_c2_443f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2335_c2_443f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2335_c2_443f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l2360_l2331_DUPLICATE_9b98 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l2360_l2331_DUPLICATE_9b98_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b93(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_443f_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_443f_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l2360_l2331_DUPLICATE_9b98_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l2360_l2331_DUPLICATE_9b98_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
