-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity ldr_0CLK_1b20325b is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldr_0CLK_1b20325b;
architecture arch of ldr_0CLK_1b20325b is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1572_c6_6937]
signal BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1572_c2_524b]
signal tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1572_c2_524b]
signal result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1572_c2_524b]
signal result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1572_c2_524b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1572_c2_524b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1572_c2_524b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1572_c2_524b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1572_c2_524b]
signal t8_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1579_c11_8f8e]
signal BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1579_c7_8a73]
signal tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1579_c7_8a73]
signal result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1579_c7_8a73]
signal result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1579_c7_8a73]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1579_c7_8a73]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1579_c7_8a73]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1579_c7_8a73]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1579_c7_8a73]
signal t8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1582_c11_b69e]
signal BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1582_c7_e9de]
signal tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1582_c7_e9de]
signal result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1582_c7_e9de]
signal result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1582_c7_e9de]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1582_c7_e9de]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1582_c7_e9de]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1582_c7_e9de]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1582_c7_e9de]
signal t8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1585_c30_b636]
signal sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1586_c22_ecf8]
signal BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_left : signed(16 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_right : signed(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_return_output : signed(17 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1588_c11_a9a4]
signal BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1588_c7_33ed]
signal tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1588_c7_33ed]
signal result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1588_c7_33ed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1588_c7_33ed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1588_c7_33ed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1588_c7_33ed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1591_c11_d2aa]
signal BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1591_c7_26a4]
signal tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1591_c7_26a4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1591_c7_26a4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1591_c7_26a4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1591_c7_26a4]
signal result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1597_c11_3738]
signal BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1597_c7_4c18]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1597_c7_4c18]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output : unsigned(0 downto 0);

function CAST_TO_int8_t_uint8_t( rhs : unsigned) return signed is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : signed(7 downto 0);

begin

      return_output := signed(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_e78e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937
BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_left,
BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_right,
BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1572_c2_524b
tmp8_MUX_uxn_opcodes_h_l1572_c2_524b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_cond,
tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue,
tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse,
tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b
result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond,
result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b
result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b
result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b
result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

-- t8_MUX_uxn_opcodes_h_l1572_c2_524b
t8_MUX_uxn_opcodes_h_l1572_c2_524b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1572_c2_524b_cond,
t8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue,
t8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse,
t8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e
BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_left,
BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_right,
BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73
tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond,
tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue,
tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse,
tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73
result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond,
result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73
result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond,
result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73
result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73
result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73
result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output);

-- t8_MUX_uxn_opcodes_h_l1579_c7_8a73
t8_MUX_uxn_opcodes_h_l1579_c7_8a73 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond,
t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue,
t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse,
t8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e
BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_left,
BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_right,
BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de
tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond,
tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue,
tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse,
tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de
result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond,
result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de
result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond,
result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de
result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de
result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de
result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output);

-- t8_MUX_uxn_opcodes_h_l1582_c7_e9de
t8_MUX_uxn_opcodes_h_l1582_c7_e9de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond,
t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue,
t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse,
t8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1585_c30_b636
sp_relative_shift_uxn_opcodes_h_l1585_c30_b636 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_ins,
sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_x,
sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_y,
sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8
BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8 : entity work.BIN_OP_PLUS_int17_t_int8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_left,
BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_right,
BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4
BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_left,
BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_right,
BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed
tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_cond,
tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue,
tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse,
tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed
result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_cond,
result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed
result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed
result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed
result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa
BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_left,
BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_right,
BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4
tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_cond,
tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue,
tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse,
tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4
result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4
result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4
result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738
BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_left,
BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_right,
BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18
result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18
result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output,
 tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
 t8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output,
 tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output,
 t8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output,
 tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output,
 t8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output,
 sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output,
 tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output,
 tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1576_c3_f774 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1580_c3_3473 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l1586_c3_56f4 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_left : signed(16 downto 0);
 variable VAR_CAST_TO_int8_t_uxn_opcodes_h_l1586_c27_0155_return_output : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_right : signed(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_return_output : signed(17 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1589_c3_2e9b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1594_c3_7415 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1582_l1572_l1579_DUPLICATE_1b39_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1572_l1591_l1588_l1582_l1579_DUPLICATE_5130_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1572_l1597_l1588_l1582_l1579_DUPLICATE_501c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1572_l1588_l1579_DUPLICATE_92d8_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1597_l1591_l1588_l1582_l1579_DUPLICATE_9c26_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1591_l1582_l1588_DUPLICATE_eba8_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1568_l1602_DUPLICATE_16b4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1594_c3_7415 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1594_c3_7415;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1576_c3_f774 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1576_c3_f774;
     VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1589_c3_2e9b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1589_c3_2e9b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1580_c3_3473 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1580_c3_3473;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_ins := VAR_ins;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_left := signed(std_logic_vector(resize(VAR_pc, 17)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse := tmp8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1591_l1582_l1588_DUPLICATE_eba8 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1591_l1582_l1588_DUPLICATE_eba8_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1582_l1572_l1579_DUPLICATE_1b39 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1582_l1572_l1579_DUPLICATE_1b39_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1579_c11_8f8e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1585_c30_b636] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_ins;
     sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_x;
     sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_return_output := sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1588_c11_a9a4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1582_c11_b69e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1597_c11_3738] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_left;
     BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_return_output := BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1597_l1591_l1588_l1582_l1579_DUPLICATE_9c26 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1597_l1591_l1588_l1582_l1579_DUPLICATE_9c26_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1572_l1588_l1579_DUPLICATE_92d8 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1572_l1588_l1579_DUPLICATE_92d8_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1572_l1597_l1588_l1582_l1579_DUPLICATE_501c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1572_l1597_l1588_l1582_l1579_DUPLICATE_501c_return_output := result.is_stack_write;

     -- CAST_TO_int8_t[uxn_opcodes_h_l1586_c27_0155] LATENCY=0
     VAR_CAST_TO_int8_t_uxn_opcodes_h_l1586_c27_0155_return_output := CAST_TO_int8_t_uint8_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1572_l1591_l1588_l1582_l1579_DUPLICATE_5130 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1572_l1591_l1588_l1582_l1579_DUPLICATE_5130_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1591_c11_d2aa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_left;
     BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output := BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1572_c6_6937] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_left;
     BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output := BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1572_c6_6937_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1579_c11_8f8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1582_c11_b69e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1588_c11_a9a4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1591_c11_d2aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1597_c11_3738_return_output;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_right := VAR_CAST_TO_int8_t_uxn_opcodes_h_l1586_c27_0155_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1572_l1588_l1579_DUPLICATE_92d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1572_l1588_l1579_DUPLICATE_92d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1572_l1588_l1579_DUPLICATE_92d8_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1582_l1572_l1579_DUPLICATE_1b39_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1582_l1572_l1579_DUPLICATE_1b39_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1582_l1572_l1579_DUPLICATE_1b39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1597_l1591_l1588_l1582_l1579_DUPLICATE_9c26_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1597_l1591_l1588_l1582_l1579_DUPLICATE_9c26_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1597_l1591_l1588_l1582_l1579_DUPLICATE_9c26_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1597_l1591_l1588_l1582_l1579_DUPLICATE_9c26_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1597_l1591_l1588_l1582_l1579_DUPLICATE_9c26_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1572_l1597_l1588_l1582_l1579_DUPLICATE_501c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1572_l1597_l1588_l1582_l1579_DUPLICATE_501c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1572_l1597_l1588_l1582_l1579_DUPLICATE_501c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1572_l1597_l1588_l1582_l1579_DUPLICATE_501c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1572_l1597_l1588_l1582_l1579_DUPLICATE_501c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1591_l1582_l1588_DUPLICATE_eba8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1591_l1582_l1588_DUPLICATE_eba8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1591_l1582_l1588_DUPLICATE_eba8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1572_l1591_l1588_l1582_l1579_DUPLICATE_5130_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1572_l1591_l1588_l1582_l1579_DUPLICATE_5130_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1572_l1591_l1588_l1582_l1579_DUPLICATE_5130_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1572_l1591_l1588_l1582_l1579_DUPLICATE_5130_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1572_l1591_l1588_l1582_l1579_DUPLICATE_5130_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1585_c30_b636_return_output;
     -- BIN_OP_PLUS[uxn_opcodes_h_l1586_c22_ecf8] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1597_c7_4c18] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1597_c7_4c18] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1591_c7_26a4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1591_c7_26a4] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_cond;
     tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output := tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1588_c7_33ed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1591_c7_26a4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;

     -- t8_MUX[uxn_opcodes_h_l1582_c7_e9de] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond <= VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond;
     t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue;
     t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output := t8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;

     -- Submodule level 2
     VAR_result_u16_value_uxn_opcodes_h_l1586_c3_56f4 := resize(unsigned(std_logic_vector(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1586_c22_ecf8_return_output)),16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1597_c7_4c18_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue := VAR_result_u16_value_uxn_opcodes_h_l1586_c3_56f4;
     -- result_u16_value_MUX[uxn_opcodes_h_l1582_c7_e9de] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output := result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1591_c7_26a4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1591_c7_26a4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1588_c7_33ed] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_cond;
     tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output := tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1588_c7_33ed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1582_c7_e9de] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;

     -- t8_MUX[uxn_opcodes_h_l1579_c7_8a73] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond <= VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond;
     t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue;
     t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output := t8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1588_c7_33ed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output := result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1591_c7_26a4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1582_c7_e9de] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;

     -- t8_MUX[uxn_opcodes_h_l1572_c2_524b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1572_c2_524b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_cond;
     t8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue;
     t8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output := t8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1582_c7_e9de] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output := result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1582_c7_e9de] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_cond;
     tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output := tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1579_c7_8a73] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1579_c7_8a73] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output := result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1588_c7_33ed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1588_c7_33ed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1588_c7_33ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1582_c7_e9de] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1579_c7_8a73] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_cond;
     tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output := tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1579_c7_8a73] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output := result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1572_c2_524b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output := result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1582_c7_e9de] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1579_c7_8a73] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1572_c2_524b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1582_c7_e9de_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1579_c7_8a73] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1579_c7_8a73] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1572_c2_524b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1572_c2_524b] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_cond;
     tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output := tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1572_c2_524b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1579_c7_8a73_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1572_c2_524b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1572_c2_524b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1568_l1602_DUPLICATE_16b4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1568_l1602_DUPLICATE_16b4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e78e(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1572_c2_524b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1572_c2_524b_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1568_l1602_DUPLICATE_16b4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e78e_uxn_opcodes_h_l1568_l1602_DUPLICATE_16b4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
