-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 41
entity lit2_0CLK_4351dde2 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit2_0CLK_4351dde2;
architecture arch of lit2_0CLK_4351dde2 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp8_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp8_high : unsigned(7 downto 0);
signal REG_COMB_tmp8_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l219_c6_361e]
signal BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l219_c2_feed]
signal tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l219_c2_feed]
signal tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(15 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l219_c2_feed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l232_c11_d2a3]
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l232_c7_fa6e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l234_c22_c57d]
signal BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l236_c11_0888]
signal BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output : unsigned(0 downto 0);

-- tmp8_high_MUX[uxn_opcodes_h_l236_c7_c7d9]
signal tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(7 downto 0);
signal tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(7 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l236_c7_c7d9]
signal tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l236_c7_c7d9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l236_c7_c7d9]
signal result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l236_c7_c7d9]
signal result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l236_c7_c7d9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l236_c7_c7d9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l236_c7_c7d9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l240_c22_869b]
signal BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l244_c11_091d]
signal BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output : unsigned(0 downto 0);

-- tmp8_low_MUX[uxn_opcodes_h_l244_c7_5e2e]
signal tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(7 downto 0);
signal tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l244_c7_5e2e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l244_c7_5e2e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l244_c7_5e2e]
signal result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l244_c7_5e2e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e393( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.u16_value := ref_toks_3;
      base.is_ram_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.is_pc_updated := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e
BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_left,
BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_right,
BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed
tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_cond,
tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed
tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_cond,
tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed
result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed
result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3
BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_left,
BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_right,
BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e
tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e
tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e
result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e
result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d
BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_left,
BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_right,
BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888
BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_left,
BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_right,
BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output);

-- tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9
tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_cond,
tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue,
tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse,
tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9
tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_cond,
tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9
result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond,
result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9
result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond,
result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b
BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_left,
BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_right,
BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d
BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_left,
BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_right,
BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output);

-- tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e
tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_cond,
tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue,
tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse,
tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e
result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_cond,
result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp8_high,
 tmp8_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output,
 tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output,
 tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l228_c3_643e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l234_c3_8a2e : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_6970 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l232_c7_fa6e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l241_c3_e90b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l240_c3_57e4 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l236_c7_c7d9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l247_c3_9c4c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_61fa_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_b286_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_57c8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_b7bb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_7a35_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l214_l252_DUPLICATE_f0e2_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp8_high : unsigned(7 downto 0);
variable REG_VAR_tmp8_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp8_high := tmp8_high;
  REG_VAR_tmp8_low := tmp8_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_right := to_unsigned(2, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_right := to_unsigned(3, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_6970 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l233_c3_6970;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_right := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l228_c3_643e := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l228_c3_643e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l247_c3_9c4c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l247_c3_9c4c;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l241_c3_e90b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l241_c3_e90b;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue := VAR_previous_ram_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue := VAR_previous_ram_read;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue := VAR_previous_ram_read;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue := VAR_previous_ram_read;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := tmp8_high;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse := tmp8_high;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue := tmp8_low;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse := tmp8_low;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_57c8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_57c8_return_output := result.is_pc_updated;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l219_c2_feed_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_61fa LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_61fa_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l219_c2_feed_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l236_c11_0888] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_left;
     BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output := BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l232_c11_d2a3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_left;
     BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output := BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_b7bb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_b7bb_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_b286 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_b286_return_output := result.u8_value;

     -- BIN_OP_PLUS[uxn_opcodes_h_l240_c22_869b] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_left;
     BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_return_output := BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l219_c6_361e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_left;
     BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output := BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l219_c2_feed_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l244_c11_091d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_left;
     BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output := BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l232_c7_fa6e_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_7a35 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_7a35_return_output := result.is_opc_done;

     -- result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l236_c7_c7d9_return_output := result.u16_value;

     -- BIN_OP_PLUS[uxn_opcodes_h_l234_c22_c57d] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_left;
     BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_return_output := BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l219_c6_361e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_d2a3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l236_c11_0888_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l244_c11_091d_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l234_c3_8a2e := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l234_c22_c57d_return_output, 16);
     VAR_result_u16_value_uxn_opcodes_h_l240_c3_57e4 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l240_c22_869b_return_output, 16);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_7a35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_7a35_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l232_l236_l244_DUPLICATE_7a35_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_57c8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l232_l244_DUPLICATE_57c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_b7bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l232_l236_DUPLICATE_b7bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_61fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_61fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_61fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_b286_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_b286_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l232_l219_l244_DUPLICATE_b286_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l219_c2_feed_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l219_c2_feed_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l219_c2_feed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l232_c7_fa6e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse := VAR_result_u16_value_FALSE_INPUT_MUX_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l236_c7_c7d9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue := VAR_result_u16_value_uxn_opcodes_h_l234_c3_8a2e;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue := VAR_result_u16_value_uxn_opcodes_h_l240_c3_57e4;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l244_c7_5e2e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output := result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l244_c7_5e2e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l244_c7_5e2e] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_cond;
     tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output := tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l244_c7_5e2e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l244_c7_5e2e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output := result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_cond;
     tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output := tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l244_c7_5e2e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_cond;
     tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output := tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output := result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l236_c7_c7d9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;
     VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_tmp8_high_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l236_c7_c7d9_return_output;
     -- tmp8_low_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l232_c7_fa6e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;

     -- tmp8_high_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_return_output := tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     REG_VAR_tmp8_high := VAR_tmp8_high_MUX_uxn_opcodes_h_l219_c2_feed_return_output;
     VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iffalse := VAR_tmp8_low_MUX_uxn_opcodes_h_l232_c7_fa6e_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- tmp8_low_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_return_output := tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l219_c2_feed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_return_output;

     -- Submodule level 5
     REG_VAR_tmp8_low := VAR_tmp8_low_MUX_uxn_opcodes_h_l219_c2_feed_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l214_l252_DUPLICATE_f0e2 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l214_l252_DUPLICATE_f0e2_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e393(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l219_c2_feed_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l219_c2_feed_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l214_l252_DUPLICATE_f0e2_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e393_uxn_opcodes_h_l214_l252_DUPLICATE_f0e2_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp8_high <= REG_VAR_tmp8_high;
REG_COMB_tmp8_low <= REG_VAR_tmp8_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp8_high <= REG_COMB_tmp8_high;
     tmp8_low <= REG_COMB_tmp8_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
