-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 52
entity add_0CLK_f62d646e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end add_0CLK_f62d646e;
architecture arch of add_0CLK_f62d646e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l854_c6_40d6]
signal BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l854_c1_34f4]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l854_c2_1a33]
signal n8_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l854_c2_1a33]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l854_c2_1a33]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l854_c2_1a33]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l854_c2_1a33]
signal result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l854_c2_1a33]
signal result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l854_c2_1a33]
signal result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l854_c2_1a33]
signal t8_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l855_c3_4913[uxn_opcodes_h_l855_c3_4913]
signal printf_uxn_opcodes_h_l855_c3_4913_uxn_opcodes_h_l855_c3_4913_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l859_c11_62d1]
signal BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l859_c7_df20]
signal n8_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l859_c7_df20]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l859_c7_df20]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l859_c7_df20]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l859_c7_df20]
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l859_c7_df20]
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l859_c7_df20]
signal result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l859_c7_df20]
signal t8_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l862_c11_a0f9]
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l862_c7_aa56]
signal n8_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l862_c7_aa56]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l862_c7_aa56]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l862_c7_aa56]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l862_c7_aa56]
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l862_c7_aa56]
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l862_c7_aa56]
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l862_c7_aa56]
signal t8_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l866_c11_8ffc]
signal BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l866_c7_d7aa]
signal n8_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l866_c7_d7aa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l866_c7_d7aa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l866_c7_d7aa]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l866_c7_d7aa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l866_c7_d7aa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l866_c7_d7aa]
signal result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l869_c11_8ca5]
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l869_c7_a2b9]
signal n8_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l869_c7_a2b9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l869_c7_a2b9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l869_c7_a2b9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l869_c7_a2b9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l869_c7_a2b9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l869_c7_a2b9]
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l872_c30_5018]
signal sp_relative_shift_uxn_opcodes_h_l872_c30_5018_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l872_c30_5018_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l872_c30_5018_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l872_c30_5018_return_output : signed(3 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l875_c21_c668]
signal BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_right : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_return_output : unsigned(8 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l877_c11_df54]
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c7_9936]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l877_c7_9936]
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l877_c7_9936]
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8cda( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6
BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_left,
BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_right,
BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_return_output);

-- n8_MUX_uxn_opcodes_h_l854_c2_1a33
n8_MUX_uxn_opcodes_h_l854_c2_1a33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l854_c2_1a33_cond,
n8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue,
n8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse,
n8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33
result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_cond,
result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

-- t8_MUX_uxn_opcodes_h_l854_c2_1a33
t8_MUX_uxn_opcodes_h_l854_c2_1a33 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l854_c2_1a33_cond,
t8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue,
t8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse,
t8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

-- printf_uxn_opcodes_h_l855_c3_4913_uxn_opcodes_h_l855_c3_4913
printf_uxn_opcodes_h_l855_c3_4913_uxn_opcodes_h_l855_c3_4913 : entity work.printf_uxn_opcodes_h_l855_c3_4913_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l855_c3_4913_uxn_opcodes_h_l855_c3_4913_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1
BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_left,
BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_right,
BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output);

-- n8_MUX_uxn_opcodes_h_l859_c7_df20
n8_MUX_uxn_opcodes_h_l859_c7_df20 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l859_c7_df20_cond,
n8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue,
n8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse,
n8_MUX_uxn_opcodes_h_l859_c7_df20_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20
result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_cond,
result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_return_output);

-- t8_MUX_uxn_opcodes_h_l859_c7_df20
t8_MUX_uxn_opcodes_h_l859_c7_df20 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l859_c7_df20_cond,
t8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue,
t8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse,
t8_MUX_uxn_opcodes_h_l859_c7_df20_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9
BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_left,
BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_right,
BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output);

-- n8_MUX_uxn_opcodes_h_l862_c7_aa56
n8_MUX_uxn_opcodes_h_l862_c7_aa56 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l862_c7_aa56_cond,
n8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue,
n8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse,
n8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56
result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_cond,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_return_output);

-- t8_MUX_uxn_opcodes_h_l862_c7_aa56
t8_MUX_uxn_opcodes_h_l862_c7_aa56 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l862_c7_aa56_cond,
t8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue,
t8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse,
t8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc
BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_left,
BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_right,
BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output);

-- n8_MUX_uxn_opcodes_h_l866_c7_d7aa
n8_MUX_uxn_opcodes_h_l866_c7_d7aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l866_c7_d7aa_cond,
n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue,
n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse,
n8_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa
result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_cond,
result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5
BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_left,
BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_right,
BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output);

-- n8_MUX_uxn_opcodes_h_l869_c7_a2b9
n8_MUX_uxn_opcodes_h_l869_c7_a2b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l869_c7_a2b9_cond,
n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue,
n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse,
n8_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9
result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_cond,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l872_c30_5018
sp_relative_shift_uxn_opcodes_h_l872_c30_5018 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l872_c30_5018_ins,
sp_relative_shift_uxn_opcodes_h_l872_c30_5018_x,
sp_relative_shift_uxn_opcodes_h_l872_c30_5018_y,
sp_relative_shift_uxn_opcodes_h_l872_c30_5018_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668
BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668 : entity work.BIN_OP_PLUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_left,
BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_right,
BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54
BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_left,
BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_right,
BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_return_output,
 n8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
 t8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output,
 n8_MUX_uxn_opcodes_h_l859_c7_df20_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_return_output,
 t8_MUX_uxn_opcodes_h_l859_c7_df20_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output,
 n8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_return_output,
 t8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output,
 n8_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output,
 n8_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output,
 sp_relative_shift_uxn_opcodes_h_l872_c30_5018_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l856_c3_73bb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l855_c3_4913_uxn_opcodes_h_l855_c3_4913_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l860_c3_bb98 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l864_c3_6b70 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_c252 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l874_c3_45b7 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l869_c7_a2b9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l875_c3_9e5b : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_return_output : unsigned(8 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_4929_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_50d4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_c10e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_3f17_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l859_l877_l869_l866_l862_DUPLICATE_701a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l883_l850_DUPLICATE_4d31_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l874_c3_45b7 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l874_c3_45b7;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_right := to_unsigned(5, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_right := to_unsigned(3, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l860_c3_bb98 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l860_c3_bb98;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_c252 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l867_c3_c252;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l864_c3_6b70 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l864_c3_6b70;
     VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l856_c3_73bb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l856_c3_73bb;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l859_c11_62d1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_left;
     BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output := BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l859_l877_l869_l866_l862_DUPLICATE_701a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l859_l877_l869_l866_l862_DUPLICATE_701a_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l872_c30_5018] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l872_c30_5018_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_ins;
     sp_relative_shift_uxn_opcodes_h_l872_c30_5018_x <= VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_x;
     sp_relative_shift_uxn_opcodes_h_l872_c30_5018_y <= VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_return_output := sp_relative_shift_uxn_opcodes_h_l872_c30_5018_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l875_c21_c668] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_left;
     BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_return_output := BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_c10e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_c10e_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_3f17 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_3f17_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_4929 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_4929_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l869_c7_a2b9] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l869_c7_a2b9_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l869_c11_8ca5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_left;
     BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output := BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l877_c11_df54] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_left;
     BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output := BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l862_c11_a0f9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_left;
     BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output := BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_50d4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_50d4_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l854_c6_40d6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_left;
     BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output := BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l866_c11_8ffc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_left;
     BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output := BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l854_c6_40d6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l859_c11_62d1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l862_c11_a0f9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l866_c11_8ffc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l869_c11_8ca5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c11_df54_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l875_c3_9e5b := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l875_c21_c668_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_4929_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_4929_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_4929_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_4929_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_4929_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l859_l877_l869_l866_l862_DUPLICATE_701a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l859_l877_l869_l866_l862_DUPLICATE_701a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l859_l877_l869_l866_l862_DUPLICATE_701a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l859_l877_l869_l866_l862_DUPLICATE_701a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l859_l877_l869_l866_l862_DUPLICATE_701a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_50d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_50d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_50d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_50d4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_50d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_c10e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_c10e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_c10e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_c10e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l859_l854_l877_l866_l862_DUPLICATE_c10e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_3f17_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_3f17_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_3f17_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_3f17_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l859_l854_l869_l866_l862_DUPLICATE_3f17_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l869_c7_a2b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l872_c30_5018_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue := VAR_result_u8_value_uxn_opcodes_h_l875_c3_9e5b;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c7_9936] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l877_c7_9936] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l869_c7_a2b9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output := result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;

     -- n8_MUX[uxn_opcodes_h_l869_c7_a2b9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l869_c7_a2b9_cond <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_cond;
     n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue;
     n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output := n8_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l877_c7_9936] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l869_c7_a2b9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;

     -- t8_MUX[uxn_opcodes_h_l862_c7_aa56] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l862_c7_aa56_cond <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_cond;
     t8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue;
     t8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output := t8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l869_c7_a2b9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l854_c1_34f4] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l855_c3_4913_uxn_opcodes_h_l855_c3_4913_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l854_c1_34f4_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse := VAR_n8_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c7_9936_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c7_9936_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c7_9936_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse := VAR_t8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l869_c7_a2b9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l866_c7_d7aa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output := result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l869_c7_a2b9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l866_c7_d7aa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l869_c7_a2b9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;

     -- n8_MUX[uxn_opcodes_h_l866_c7_d7aa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l866_c7_d7aa_cond <= VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_cond;
     n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue;
     n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output := n8_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;

     -- t8_MUX[uxn_opcodes_h_l859_c7_df20] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l859_c7_df20_cond <= VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_cond;
     t8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue;
     t8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_return_output := t8_MUX_uxn_opcodes_h_l859_c7_df20_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l866_c7_d7aa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;

     -- printf_uxn_opcodes_h_l855_c3_4913[uxn_opcodes_h_l855_c3_4913] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l855_c3_4913_uxn_opcodes_h_l855_c3_4913_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l855_c3_4913_uxn_opcodes_h_l855_c3_4913_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse := VAR_n8_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l869_c7_a2b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse := VAR_t8_MUX_uxn_opcodes_h_l859_c7_df20_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l866_c7_d7aa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l866_c7_d7aa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l862_c7_aa56] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;

     -- n8_MUX[uxn_opcodes_h_l862_c7_aa56] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l862_c7_aa56_cond <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_cond;
     n8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue;
     n8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output := n8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;

     -- t8_MUX[uxn_opcodes_h_l854_c2_1a33] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l854_c2_1a33_cond <= VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_cond;
     t8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue;
     t8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output := t8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l866_c7_d7aa] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l862_c7_aa56] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_cond;
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_return_output := result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l862_c7_aa56] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse := VAR_n8_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l866_c7_d7aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;
     -- n8_MUX[uxn_opcodes_h_l859_c7_df20] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l859_c7_df20_cond <= VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_cond;
     n8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_iftrue;
     n8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_return_output := n8_MUX_uxn_opcodes_h_l859_c7_df20_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l859_c7_df20] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l862_c7_aa56] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l862_c7_aa56] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l862_c7_aa56] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l859_c7_df20] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_cond;
     result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_return_output := result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l859_c7_df20] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse := VAR_n8_MUX_uxn_opcodes_h_l859_c7_df20_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l862_c7_aa56_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l859_c7_df20_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l859_c7_df20_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l859_c7_df20] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l854_c2_1a33] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_cond;
     result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_return_output := result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l859_c7_df20] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l859_c7_df20] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output;

     -- n8_MUX[uxn_opcodes_h_l854_c2_1a33] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l854_c2_1a33_cond <= VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_cond;
     n8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue;
     n8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output := n8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l854_c2_1a33] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l854_c2_1a33] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l859_c7_df20_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l859_c7_df20_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l859_c7_df20_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l854_c2_1a33] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l854_c2_1a33] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l854_c2_1a33] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l883_l850_DUPLICATE_4d31 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l883_l850_DUPLICATE_4d31_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8cda(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l854_c2_1a33_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l854_c2_1a33_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l883_l850_DUPLICATE_4d31_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8cda_uxn_opcodes_h_l883_l850_DUPLICATE_4d31_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
