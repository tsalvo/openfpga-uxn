-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity neq2_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end neq2_0CLK_85d5529e;
architecture arch of neq2_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1162_c6_d538]
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal n16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1162_c2_b7db]
signal t16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1170_c11_2c20]
signal BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1170_c7_f501]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1170_c7_f501]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1170_c7_f501]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1170_c7_f501]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1170_c7_f501]
signal result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1170_c7_f501]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1170_c7_f501]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1170_c7_f501]
signal n16_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1170_c7_f501]
signal t16_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1173_c11_1452]
signal BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(0 downto 0);

-- n16_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal n16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l1173_c7_ceac]
signal t16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1177_c30_677e]
signal sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1179_c11_480f]
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1179_c7_c6c4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1179_c7_c6c4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1179_c7_c6c4]
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1179_c7_c6c4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1179_c7_c6c4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(3 downto 0);

-- n16_MUX[uxn_opcodes_h_l1179_c7_c6c4]
signal n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
signal n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(15 downto 0);
signal n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1184_c21_7bb2]
signal BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_left : unsigned(15 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_right : unsigned(15 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1184_c21_a49f]
signal MUX_uxn_opcodes_h_l1184_c21_a49f_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1184_c21_a49f_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1184_c21_a49f_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1184_c21_a49f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1186_c11_527d]
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1186_c7_e0e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1186_c7_e0e5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_stack_operation_16bit := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_stack_write := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_left,
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_right,
BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db
result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- n16_MUX_uxn_opcodes_h_l1162_c2_b7db
n16_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
n16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- t16_MUX_uxn_opcodes_h_l1162_c2_b7db
t16_MUX_uxn_opcodes_h_l1162_c2_b7db : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond,
t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue,
t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse,
t16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20
BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_left,
BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_right,
BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501
result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501
result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501
result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501
result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501
result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- n16_MUX_uxn_opcodes_h_l1170_c7_f501
n16_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
n16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
n16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
n16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- t16_MUX_uxn_opcodes_h_l1170_c7_f501
t16_MUX_uxn_opcodes_h_l1170_c7_f501 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1170_c7_f501_cond,
t16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue,
t16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse,
t16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452
BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_left,
BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_right,
BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac
result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac
result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac
result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac
result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac
result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- n16_MUX_uxn_opcodes_h_l1173_c7_ceac
n16_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
n16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- t16_MUX_uxn_opcodes_h_l1173_c7_ceac
t16_MUX_uxn_opcodes_h_l1173_c7_ceac : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond,
t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue,
t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse,
t16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1177_c30_677e
sp_relative_shift_uxn_opcodes_h_l1177_c30_677e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_ins,
sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_x,
sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_y,
sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_left,
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_right,
BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4
result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output);

-- n16_MUX_uxn_opcodes_h_l1179_c7_c6c4
n16_MUX_uxn_opcodes_h_l1179_c7_c6c4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond,
n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue,
n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse,
n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2
BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2 : entity work.BIN_OP_EQ_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_left,
BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_right,
BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_return_output);

-- MUX_uxn_opcodes_h_l1184_c21_a49f
MUX_uxn_opcodes_h_l1184_c21_a49f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1184_c21_a49f_cond,
MUX_uxn_opcodes_h_l1184_c21_a49f_iftrue,
MUX_uxn_opcodes_h_l1184_c21_a49f_iffalse,
MUX_uxn_opcodes_h_l1184_c21_a49f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d
BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_left,
BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_right,
BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5
result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5
result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 n16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 t16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 n16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 t16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 n16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 t16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output,
 sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output,
 n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_return_output,
 MUX_uxn_opcodes_h_l1184_c21_a49f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1167_c3_74e6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1171_c3_72c5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1183_c3_ae9a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse : unsigned(15 downto 0);
 variable VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1170_l1162_l1179_DUPLICATE_67e6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1173_l1170_l1162_l1179_DUPLICATE_d5e0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1173_l1170_l1162_DUPLICATE_d1b5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1162_DUPLICATE_9ee2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1173_l1170_DUPLICATE_1064_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1179_DUPLICATE_ff86_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1173_l1179_DUPLICATE_58f6_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1158_l1191_DUPLICATE_1692_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n16 := n16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_y := resize(to_signed(-3, 3), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1171_c3_72c5 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1171_c3_72c5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1167_c3_74e6 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1167_c3_74e6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1183_c3_ae9a := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1183_c3_ae9a;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_ins := VAR_ins;
     VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := n16;
     VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse := n16;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_left := VAR_previous_stack_read;
     VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_right := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1162_DUPLICATE_9ee2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1162_DUPLICATE_9ee2_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1173_l1170_DUPLICATE_1064 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1173_l1170_DUPLICATE_1064_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1173_l1170_l1162_DUPLICATE_d1b5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1173_l1170_l1162_DUPLICATE_d1b5_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1162_c6_d538] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_left;
     BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output := BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1170_c11_2c20] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_left;
     BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output := BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1186_c11_527d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1177_c30_677e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_ins;
     sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_x;
     sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_return_output := sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1173_l1179_DUPLICATE_58f6 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1173_l1179_DUPLICATE_58f6_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1170_l1162_l1179_DUPLICATE_67e6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1170_l1162_l1179_DUPLICATE_67e6_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1179_DUPLICATE_ff86 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1179_DUPLICATE_ff86_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1184_c21_7bb2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1179_c11_480f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1173_l1170_l1162_l1179_DUPLICATE_d5e0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1173_l1170_l1162_l1179_DUPLICATE_d5e0_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1173_c11_1452] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_left;
     BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output := BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;

     -- Submodule level 1
     VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1162_c6_d538_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1170_c11_2c20_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1173_c11_1452_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1179_c11_480f_return_output;
     VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1184_c21_7bb2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1186_c11_527d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1173_l1170_l1162_DUPLICATE_d1b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1173_l1170_l1162_DUPLICATE_d1b5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1173_l1170_l1162_DUPLICATE_d1b5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1179_DUPLICATE_ff86_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1179_DUPLICATE_ff86_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1179_DUPLICATE_ff86_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1179_DUPLICATE_ff86_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1170_l1162_l1179_DUPLICATE_67e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1170_l1162_l1179_DUPLICATE_67e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1170_l1162_l1179_DUPLICATE_67e6_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1173_l1170_DUPLICATE_1064_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l1173_l1170_DUPLICATE_1064_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1162_DUPLICATE_9ee2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1162_DUPLICATE_9ee2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1162_DUPLICATE_9ee2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1173_l1170_l1186_l1162_DUPLICATE_9ee2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1173_l1179_DUPLICATE_58f6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1173_l1179_DUPLICATE_58f6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1173_l1170_l1162_l1179_DUPLICATE_d5e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1173_l1170_l1162_l1179_DUPLICATE_d5e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1173_l1170_l1162_l1179_DUPLICATE_d5e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1173_l1170_l1162_l1179_DUPLICATE_d5e0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1177_c30_677e_return_output;
     -- n16_MUX[uxn_opcodes_h_l1179_c7_c6c4] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond <= VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond;
     n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue;
     n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output := n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1186_c7_e0e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output;

     -- MUX[uxn_opcodes_h_l1184_c21_a49f] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1184_c21_a49f_cond <= VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_cond;
     MUX_uxn_opcodes_h_l1184_c21_a49f_iftrue <= VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_iftrue;
     MUX_uxn_opcodes_h_l1184_c21_a49f_iffalse <= VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_return_output := MUX_uxn_opcodes_h_l1184_c21_a49f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1186_c7_e0e5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1179_c7_c6c4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1179_c7_c6c4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;

     -- t16_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := t16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue := VAR_MUX_uxn_opcodes_h_l1184_c21_a49f_return_output;
     VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1186_c7_e0e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- t16_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     t16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     t16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := t16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1179_c7_c6c4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1179_c7_c6c4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- n16_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := n16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1179_c7_c6c4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;

     -- Submodule level 3
     VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1179_c7_c6c4_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_t16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- t16_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := t16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- n16_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     n16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     n16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := n16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1173_c7_ceac] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output := result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;

     -- Submodule level 4
     VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_n16_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1173_c7_ceac_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- n16_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     n16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := n16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1170_c7_f501] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- Submodule level 5
     REG_VAR_n16 := VAR_n16_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1170_c7_f501_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1162_c2_b7db] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1158_l1191_DUPLICATE_1692 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1158_l1191_DUPLICATE_1692_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1162_c2_b7db_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1158_l1191_DUPLICATE_1692_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9d9a_uxn_opcodes_h_l1158_l1191_DUPLICATE_1692_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n16 <= REG_VAR_n16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n16 <= REG_COMB_n16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
