-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity mul_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end mul_0CLK_64d180f1;
architecture arch of mul_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1969_c6_2a41]
signal BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1969_c2_ab8b]
signal t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1982_c11_6d88]
signal BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1982_c7_0320]
signal n8_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1982_c7_0320]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1982_c7_0320]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1982_c7_0320]
signal result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1982_c7_0320]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1982_c7_0320]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1982_c7_0320]
signal t8_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1985_c11_c25c]
signal BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1985_c7_9606]
signal n8_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1985_c7_9606]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1985_c7_9606]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1985_c7_9606]
signal result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1985_c7_9606]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1985_c7_9606]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1985_c7_9606]
signal t8_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1988_c11_eb1c]
signal BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1988_c7_e058]
signal n8_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1988_c7_e058]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1988_c7_e058]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1988_c7_e058]
signal result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1988_c7_e058]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1988_c7_e058]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1990_c30_cdab]
signal sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_return_output : signed(3 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1993_c21_c815]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_return_output : unsigned(15 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8b52( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_ram_write := ref_toks_7;
      base.is_vram_write := ref_toks_8;
      base.u8_value := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41
BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_left,
BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_right,
BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output);

-- n8_MUX_uxn_opcodes_h_l1969_c2_ab8b
n8_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- t8_MUX_uxn_opcodes_h_l1969_c2_ab8b
t8_MUX_uxn_opcodes_h_l1969_c2_ab8b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond,
t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue,
t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse,
t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88
BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_left,
BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_right,
BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output);

-- n8_MUX_uxn_opcodes_h_l1982_c7_0320
n8_MUX_uxn_opcodes_h_l1982_c7_0320 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1982_c7_0320_cond,
n8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue,
n8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse,
n8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_cond,
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_return_output);

-- t8_MUX_uxn_opcodes_h_l1982_c7_0320
t8_MUX_uxn_opcodes_h_l1982_c7_0320 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1982_c7_0320_cond,
t8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue,
t8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse,
t8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c
BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_left,
BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_right,
BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output);

-- n8_MUX_uxn_opcodes_h_l1985_c7_9606
n8_MUX_uxn_opcodes_h_l1985_c7_9606 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1985_c7_9606_cond,
n8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue,
n8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse,
n8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_cond,
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_return_output);

-- t8_MUX_uxn_opcodes_h_l1985_c7_9606
t8_MUX_uxn_opcodes_h_l1985_c7_9606 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1985_c7_9606_cond,
t8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue,
t8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse,
t8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c
BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_left,
BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_right,
BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output);

-- n8_MUX_uxn_opcodes_h_l1988_c7_e058
n8_MUX_uxn_opcodes_h_l1988_c7_e058 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1988_c7_e058_cond,
n8_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue,
n8_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse,
n8_MUX_uxn_opcodes_h_l1988_c7_e058_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_cond,
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab
sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_ins,
sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_x,
sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_y,
sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815 : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output,
 n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output,
 n8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_return_output,
 t8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output,
 n8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_return_output,
 t8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output,
 n8_MUX_uxn_opcodes_h_l1988_c7_e058_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_return_output,
 sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1974_c3_495b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1979_c3_1346 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1983_c3_df5b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_uxn_opcodes_h_l1993_c3_fd3e : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1992_c3_2fdf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1982_l1985_l1969_l1988_DUPLICATE_4982_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b40b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b072_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_2f97_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_7a59_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1997_l1965_DUPLICATE_24b0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1974_c3_495b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1974_c3_495b;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1992_c3_2fdf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1992_c3_2fdf;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1983_c3_df5b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1983_c3_df5b;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_right := to_unsigned(3, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1979_c3_1346 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1979_c3_1346;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_left := VAR_phase;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_2f97 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_2f97_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b072 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b072_return_output := result.is_stack_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1988_c11_eb1c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1985_c11_c25c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_7a59 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_7a59_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1990_c30_cdab] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_ins;
     sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_x;
     sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_return_output := sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1982_c11_6d88] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_left;
     BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output := BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1969_c6_2a41] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_left;
     BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output := BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output := result.is_pc_updated;

     -- BIN_OP_INFERRED_MULT[uxn_opcodes_h_l1993_c21_c815] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b40b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b40b_return_output := result.sp_relative_shift;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1982_l1985_l1969_l1988_DUPLICATE_4982 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1982_l1985_l1969_l1988_DUPLICATE_4982_return_output := result.u8_value;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1969_c6_2a41_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1982_c11_6d88_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1985_c11_c25c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1988_c11_eb1c_return_output;
     VAR_result_u8_value_uxn_opcodes_h_l1993_c3_fd3e := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_h_l1993_c21_c815_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b40b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b40b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b40b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_2f97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_2f97_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_2f97_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b072_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b072_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1982_l1985_l1988_DUPLICATE_b072_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_7a59_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1985_l1988_DUPLICATE_7a59_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1982_l1985_l1969_l1988_DUPLICATE_4982_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1982_l1985_l1969_l1988_DUPLICATE_4982_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1982_l1985_l1969_l1988_DUPLICATE_4982_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1982_l1985_l1969_l1988_DUPLICATE_4982_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1969_c2_ab8b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1990_c30_cdab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue := VAR_result_u8_value_uxn_opcodes_h_l1993_c3_fd3e;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1988_c7_e058] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1988_c7_e058] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_return_output := result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1988_c7_e058] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1988_c7_e058] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;

     -- t8_MUX[uxn_opcodes_h_l1985_c7_9606] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1985_c7_9606_cond <= VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_cond;
     t8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue;
     t8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output := t8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1988_c7_e058] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1988_c7_e058_cond <= VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_cond;
     n8_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue;
     n8_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_return_output := n8_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1988_c7_e058] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1988_c7_e058_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1985_c7_9606] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1985_c7_9606] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;

     -- t8_MUX[uxn_opcodes_h_l1982_c7_0320] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1982_c7_0320_cond <= VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_cond;
     t8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue;
     t8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output := t8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1985_c7_9606] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_return_output := result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;

     -- n8_MUX[uxn_opcodes_h_l1985_c7_9606] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1985_c7_9606_cond <= VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_cond;
     n8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue;
     n8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output := n8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1985_c7_9606] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1985_c7_9606] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1985_c7_9606_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1982_c7_0320] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1982_c7_0320] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;

     -- n8_MUX[uxn_opcodes_h_l1982_c7_0320] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1982_c7_0320_cond <= VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_cond;
     n8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue;
     n8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output := n8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;

     -- t8_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1982_c7_0320] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1982_c7_0320] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_return_output := result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1982_c7_0320] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1982_c7_0320_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1969_c2_ab8b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_cond;
     n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iftrue;
     n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output := n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1997_l1965_DUPLICATE_24b0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1997_l1965_DUPLICATE_24b0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8b52(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1969_c2_ab8b_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1997_l1965_DUPLICATE_24b0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8b52_uxn_opcodes_h_l1997_l1965_DUPLICATE_24b0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
