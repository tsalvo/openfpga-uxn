-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity lit2_0CLK_edc09f97 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit2_0CLK_edc09f97;
architecture arch of lit2_0CLK_edc09f97 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l214_c6_4a7c]
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l214_c1_f658]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l214_c2_bac2]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l214_c2_bac2]
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l214_c2_bac2]
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l214_c2_bac2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l214_c2_bac2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l214_c2_bac2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l214_c2_bac2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l214_c2_bac2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(3 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l214_c2_bac2]
signal tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l215_c3_f560[uxn_opcodes_h_l215_c3_f560]
signal printf_uxn_opcodes_h_l215_c3_f560_uxn_opcodes_h_l215_c3_f560_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l221_c11_44ab]
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l221_c7_a6f4]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l221_c7_a6f4]
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l221_c7_a6f4]
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l221_c7_a6f4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l221_c7_a6f4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l221_c7_a6f4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l221_c7_a6f4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(3 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l221_c7_a6f4]
signal tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l223_c22_2421]
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l225_c11_1037]
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l225_c7_b750]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l225_c7_b750]
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l225_c7_b750]
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l225_c7_b750]
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l225_c7_b750]
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l225_c7_b750]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(3 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l225_c7_b750]
signal tmp16_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l227_c3_f747]
signal CONST_SL_8_uxn_opcodes_h_l227_c3_f747_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l227_c3_f747_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l229_c11_24fa]
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l229_c7_6342]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l229_c7_6342]
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(15 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l229_c7_6342]
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l229_c7_6342]
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l229_c7_6342]
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l229_c7_6342]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(3 downto 0);

-- tmp16_MUX[uxn_opcodes_h_l229_c7_6342]
signal tmp16_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(15 downto 0);
signal tmp16_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l230_c3_84d4]
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_return_output : unsigned(15 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l232_c22_3730]
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_right : unsigned(1 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l237_c11_accb]
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l237_c7_8969]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l237_c7_8969]
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l237_c7_8969]
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l237_c7_8969]
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l237_c7_8969]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(3 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l240_c31_f124]
signal CONST_SR_8_uxn_opcodes_h_l240_c31_f124_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l240_c31_f124_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l242_c11_0d46]
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l242_c7_e762]
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l242_c7_e762]
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_2af2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_pc_updated := ref_toks_1;
      base.u16_value := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.is_opc_done := ref_toks_6;
      base.is_stack_write := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c
BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_left,
BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_right,
BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2
result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2
result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- tmp16_MUX_uxn_opcodes_h_l214_c2_bac2
tmp16_MUX_uxn_opcodes_h_l214_c2_bac2 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_cond,
tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue,
tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse,
tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

-- printf_uxn_opcodes_h_l215_c3_f560_uxn_opcodes_h_l215_c3_f560
printf_uxn_opcodes_h_l215_c3_f560_uxn_opcodes_h_l215_c3_f560 : entity work.printf_uxn_opcodes_h_l215_c3_f560_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l215_c3_f560_uxn_opcodes_h_l215_c3_f560_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab
BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_left,
BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_right,
BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4
result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4
result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output);

-- tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4
tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_cond,
tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue,
tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse,
tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_left,
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_right,
BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037
BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_left,
BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_right,
BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_cond,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_cond,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_return_output);

-- tmp16_MUX_uxn_opcodes_h_l225_c7_b750
tmp16_MUX_uxn_opcodes_h_l225_c7_b750 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l225_c7_b750_cond,
tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iftrue,
tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iffalse,
tmp16_MUX_uxn_opcodes_h_l225_c7_b750_return_output);

-- CONST_SL_8_uxn_opcodes_h_l227_c3_f747
CONST_SL_8_uxn_opcodes_h_l227_c3_f747 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l227_c3_f747_x,
CONST_SL_8_uxn_opcodes_h_l227_c3_f747_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa
BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_left,
BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_right,
BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342
result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_cond,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342
result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_cond,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_return_output);

-- tmp16_MUX_uxn_opcodes_h_l229_c7_6342
tmp16_MUX_uxn_opcodes_h_l229_c7_6342 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
tmp16_MUX_uxn_opcodes_h_l229_c7_6342_cond,
tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iftrue,
tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iffalse,
tmp16_MUX_uxn_opcodes_h_l229_c7_6342_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4
BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4 : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_left,
BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_right,
BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730 : entity work.BIN_OP_PLUS_uint16_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_left,
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_right,
BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb
BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_left,
BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_right,
BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_cond,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_return_output);

-- CONST_SR_8_uxn_opcodes_h_l240_c31_f124
CONST_SR_8_uxn_opcodes_h_l240_c31_f124 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l240_c31_f124_x,
CONST_SR_8_uxn_opcodes_h_l240_c31_f124_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46
BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_left,
BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_right,
BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output,
 tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_return_output,
 tmp16_MUX_uxn_opcodes_h_l225_c7_b750_return_output,
 CONST_SL_8_uxn_opcodes_h_l227_c3_f747_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_return_output,
 tmp16_MUX_uxn_opcodes_h_l229_c7_6342_return_output,
 BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_return_output,
 CONST_SR_8_uxn_opcodes_h_l240_c31_f124_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_cce0 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_bac2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l215_c3_f560_uxn_opcodes_h_l215_c3_f560_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l223_c3_a586 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_a6f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_return_output : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_f747_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_f747_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_uxn_opcodes_h_l232_c3_ae88 : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_bf02 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iftrue : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iffalse : unsigned(15 downto 0);
 variable VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_return_output : unsigned(16 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_8c30_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_8e13 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_f124_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_f124_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_9a30_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_b770_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_dfe8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l221_l242_l225_l237_DUPLICATE_a282_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_5184_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l221_l242_l229_l225_l237_DUPLICATE_9235_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l230_l226_DUPLICATE_79e6_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_c414_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2af2_uxn_opcodes_h_l247_l209_DUPLICATE_ae0e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp16 := tmp16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_bf02 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l234_c3_bf02;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_cce0 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l217_c3_cce0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_right := to_unsigned(5, 3);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_8e13 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l239_c3_8e13;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_right := to_unsigned(3, 2);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_right := to_unsigned(4, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_left := VAR_pc;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_left := VAR_pc;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_left := tmp16;
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_f124_x := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue := tmp16;
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iffalse := tmp16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_b770 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_b770_return_output := result.is_pc_updated;

     -- result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_a6f4_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_c414 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_c414_return_output := result.u16_value;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l230_l226_DUPLICATE_79e6 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l230_l226_DUPLICATE_79e6_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_ram_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l221_l242_l229_l225_l237_DUPLICATE_9235 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l221_l242_l229_l225_l237_DUPLICATE_9235_return_output := result.is_opc_done;

     -- CONST_SR_8[uxn_opcodes_h_l240_c31_f124] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l240_c31_f124_x <= VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_f124_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_f124_return_output := CONST_SR_8_uxn_opcodes_h_l240_c31_f124_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l221_c11_44ab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_left;
     BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output := BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l214_c6_4a7c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_left;
     BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output := BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l237_c11_accb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_left;
     BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output := BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l223_c22_2421] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_left;
     BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_return_output := BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_return_output;

     -- BIN_OP_PLUS[uxn_opcodes_h_l232_c22_3730] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_left;
     BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_return_output := BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_bac2_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_dfe8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_dfe8_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l229_c11_24fa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_left;
     BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output := BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_5184 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_5184_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l242_c11_0d46] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_left;
     BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_return_output := BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l221_l242_l225_l237_DUPLICATE_a282 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l221_l242_l225_l237_DUPLICATE_a282_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l225_c11_1037] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_left;
     BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output := BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l214_c6_4a7c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l221_c11_44ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l225_c11_1037_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l229_c11_24fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l237_c11_accb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l242_c11_0d46_return_output;
     VAR_result_u16_value_uxn_opcodes_h_l223_c3_a586 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l223_c22_2421_return_output, 16);
     VAR_result_u16_value_uxn_opcodes_h_l232_c3_ae88 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l232_c22_3730_return_output, 16);
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l230_l226_DUPLICATE_79e6_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_f747_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l230_l226_DUPLICATE_79e6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_c414_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l229_l225_DUPLICATE_c414_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l221_l242_l229_l225_l237_DUPLICATE_9235_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l221_l242_l229_l225_l237_DUPLICATE_9235_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l221_l242_l229_l225_l237_DUPLICATE_9235_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l221_l242_l229_l225_l237_DUPLICATE_9235_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l221_l242_l229_l225_l237_DUPLICATE_9235_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_b770_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_b770_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_b770_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_b770_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l221_l242_l225_l237_DUPLICATE_a282_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l221_l242_l225_l237_DUPLICATE_a282_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l221_l242_l225_l237_DUPLICATE_a282_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l221_l242_l225_l237_DUPLICATE_a282_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l214_l221_l242_l225_l237_DUPLICATE_a282_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_5184_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_5184_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_5184_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_5184_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_dfe8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_dfe8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_dfe8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l214_l221_l225_l237_DUPLICATE_dfe8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse := VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l221_c7_a6f4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l214_c2_bac2_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue := VAR_result_u16_value_uxn_opcodes_h_l223_c3_a586;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue := VAR_result_u16_value_uxn_opcodes_h_l232_c3_ae88;
     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l214_c1_f658] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l242_c7_e762] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l229_c7_6342] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_cond;
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output := result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l242_c7_e762] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l237_c7_8969] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l227_c3_f747] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l227_c3_f747_x <= VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_f747_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_f747_return_output := CONST_SL_8_uxn_opcodes_h_l227_c3_f747_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l237_c7_8969] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l230_c3_84d4] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_left;
     BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_return_output := BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l240_c21_9a30] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_9a30_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l240_c31_f124_return_output);

     -- Submodule level 2
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l240_c21_9a30_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l227_c3_f747_return_output;
     VAR_printf_uxn_opcodes_h_l215_c3_f560_uxn_opcodes_h_l215_c3_f560_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l214_c1_f658_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l242_c7_e762_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l237_c7_8969_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l242_c7_e762_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l237_c7_8969_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l229_c7_6342] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l237_c7_8969] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l229_c7_6342] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l225_c7_b750] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_cond;
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output := result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l235_c21_8c30] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_8c30_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l230_c3_84d4_return_output);

     -- tmp16_MUX[uxn_opcodes_h_l229_c7_6342] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l229_c7_6342_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_cond;
     tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iftrue;
     tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_return_output := tmp16_MUX_uxn_opcodes_h_l229_c7_6342_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l237_c7_8969] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l237_c7_8969] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_cond;
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_return_output := result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_return_output;

     -- printf_uxn_opcodes_h_l215_c3_f560[uxn_opcodes_h_l215_c3_f560] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l215_c3_f560_uxn_opcodes_h_l215_c3_f560_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l215_c3_f560_uxn_opcodes_h_l215_c3_f560_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l235_c21_8c30_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l237_c7_8969_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l229_c7_6342_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l237_c7_8969_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l229_c7_6342_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l237_c7_8969_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l229_c7_6342_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond;
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output := result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l229_c7_6342] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l229_c7_6342] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_cond;
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output := result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l229_c7_6342] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l225_c7_b750] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l225_c7_b750] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_return_output;

     -- tmp16_MUX[uxn_opcodes_h_l225_c7_b750] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l225_c7_b750_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_cond;
     tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iftrue;
     tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_return_output := tmp16_MUX_uxn_opcodes_h_l225_c7_b750_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l229_c7_6342_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l225_c7_b750_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l229_c7_6342_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l225_c7_b750_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l229_c7_6342_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l225_c7_b750_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_cond;
     tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue;
     tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output := tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l225_c7_b750] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_cond;
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output := result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l225_c7_b750] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l225_c7_b750] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l225_c7_b750_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l225_c7_b750_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l225_c7_b750_return_output;
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_tmp16_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;
     -- tmp16_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output := result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l221_c7_a6f4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l221_c7_a6f4_return_output;
     REG_VAR_tmp16 := VAR_tmp16_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l214_c2_bac2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output := result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_2af2_uxn_opcodes_h_l247_l209_DUPLICATE_ae0e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2af2_uxn_opcodes_h_l247_l209_DUPLICATE_ae0e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_2af2(
     result,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l214_c2_bac2_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l214_c2_bac2_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2af2_uxn_opcodes_h_l247_l209_DUPLICATE_ae0e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2af2_uxn_opcodes_h_l247_l209_DUPLICATE_ae0e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp16 <= REG_VAR_tmp16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp16 <= REG_COMB_tmp16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
