-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity and_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_64d180f1;
architecture arch of and_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l904_c6_72b8]
signal BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l904_c2_d47e]
signal n8_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l904_c2_d47e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l904_c2_d47e]
signal t8_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l917_c11_9d7b]
signal BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l917_c7_722f]
signal n8_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l917_c7_722f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l917_c7_722f]
signal result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l917_c7_722f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l917_c7_722f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l917_c7_722f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l917_c7_722f]
signal t8_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l920_c11_db82]
signal BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l920_c7_94ca]
signal n8_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l920_c7_94ca]
signal result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l920_c7_94ca]
signal result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l920_c7_94ca]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l920_c7_94ca]
signal result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l920_c7_94ca]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l920_c7_94ca]
signal t8_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l923_c11_bbc8]
signal BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l923_c7_0425]
signal n8_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l923_c7_0425]
signal result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l923_c7_0425]
signal result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l923_c7_0425]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l923_c7_0425]
signal result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l923_c7_0425]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l925_c30_66df]
signal sp_relative_shift_uxn_opcodes_h_l925_c30_66df_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l925_c30_66df_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l925_c30_66df_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l925_c30_66df_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l928_c21_d6fa]
signal BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8
BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_left,
BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_right,
BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output);

-- n8_MUX_uxn_opcodes_h_l904_c2_d47e
n8_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
n8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
n8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
n8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e
result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e
result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e
result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e
result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e
result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e
result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e
result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- t8_MUX_uxn_opcodes_h_l904_c2_d47e
t8_MUX_uxn_opcodes_h_l904_c2_d47e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l904_c2_d47e_cond,
t8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue,
t8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse,
t8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b
BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_left,
BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_right,
BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output);

-- n8_MUX_uxn_opcodes_h_l917_c7_722f
n8_MUX_uxn_opcodes_h_l917_c7_722f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l917_c7_722f_cond,
n8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue,
n8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse,
n8_MUX_uxn_opcodes_h_l917_c7_722f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f
result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f
result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_cond,
result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f
result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f
result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_return_output);

-- t8_MUX_uxn_opcodes_h_l917_c7_722f
t8_MUX_uxn_opcodes_h_l917_c7_722f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l917_c7_722f_cond,
t8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue,
t8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse,
t8_MUX_uxn_opcodes_h_l917_c7_722f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82
BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_left,
BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_right,
BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output);

-- n8_MUX_uxn_opcodes_h_l920_c7_94ca
n8_MUX_uxn_opcodes_h_l920_c7_94ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l920_c7_94ca_cond,
n8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue,
n8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse,
n8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca
result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca
result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_cond,
result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca
result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca
result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_return_output);

-- t8_MUX_uxn_opcodes_h_l920_c7_94ca
t8_MUX_uxn_opcodes_h_l920_c7_94ca : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l920_c7_94ca_cond,
t8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue,
t8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse,
t8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8
BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_left,
BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_right,
BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output);

-- n8_MUX_uxn_opcodes_h_l923_c7_0425
n8_MUX_uxn_opcodes_h_l923_c7_0425 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l923_c7_0425_cond,
n8_MUX_uxn_opcodes_h_l923_c7_0425_iftrue,
n8_MUX_uxn_opcodes_h_l923_c7_0425_iffalse,
n8_MUX_uxn_opcodes_h_l923_c7_0425_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425
result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425
result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_cond,
result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425
result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425
result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_return_output);

-- sp_relative_shift_uxn_opcodes_h_l925_c30_66df
sp_relative_shift_uxn_opcodes_h_l925_c30_66df : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l925_c30_66df_ins,
sp_relative_shift_uxn_opcodes_h_l925_c30_66df_x,
sp_relative_shift_uxn_opcodes_h_l925_c30_66df_y,
sp_relative_shift_uxn_opcodes_h_l925_c30_66df_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa
BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_left,
BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_right,
BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output,
 n8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 t8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output,
 n8_MUX_uxn_opcodes_h_l917_c7_722f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_return_output,
 t8_MUX_uxn_opcodes_h_l917_c7_722f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output,
 n8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_return_output,
 t8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output,
 n8_MUX_uxn_opcodes_h_l923_c7_0425_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_return_output,
 sp_relative_shift_uxn_opcodes_h_l925_c30_66df_return_output,
 BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l909_c3_ea80 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l914_c3_fc26 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l918_c3_aaef : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l927_c3_3fdc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l920_l904_l923_l917_DUPLICATE_74fb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_edf3_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_1bef_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_ce8c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l920_l923_DUPLICATE_fe23_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l932_l900_DUPLICATE_eb2d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l927_c3_3fdc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l927_c3_3fdc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l914_c3_fc26 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l914_c3_fc26;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l918_c3_aaef := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l918_c3_aaef;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l909_c3_ea80 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l909_c3_ea80;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_right := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse := t8;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l920_l923_DUPLICATE_fe23 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l920_l923_DUPLICATE_fe23_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l904_c2_d47e_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l920_c11_db82] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_left;
     BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output := BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l923_c11_bbc8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_left;
     BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output := BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l928_c21_d6fa] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_left;
     BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_return_output := BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l920_l904_l923_l917_DUPLICATE_74fb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l920_l904_l923_l917_DUPLICATE_74fb_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_edf3 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_edf3_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_ce8c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_ce8c_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l917_c11_9d7b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_left;
     BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output := BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l904_c2_d47e_return_output := result.is_ram_write;

     -- sp_relative_shift[uxn_opcodes_h_l925_c30_66df] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l925_c30_66df_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_ins;
     sp_relative_shift_uxn_opcodes_h_l925_c30_66df_x <= VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_x;
     sp_relative_shift_uxn_opcodes_h_l925_c30_66df_y <= VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_return_output := sp_relative_shift_uxn_opcodes_h_l925_c30_66df_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l904_c2_d47e_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l904_c6_72b8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_left;
     BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output := BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l904_c2_d47e_return_output := result.is_vram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_1bef LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_1bef_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l928_c21_d6fa_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l904_c6_72b8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l917_c11_9d7b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l920_c11_db82_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l923_c11_bbc8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_1bef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_1bef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_1bef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_ce8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_ce8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_ce8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_edf3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_edf3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l920_l923_l917_DUPLICATE_edf3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l920_l923_DUPLICATE_fe23_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l920_l923_DUPLICATE_fe23_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l920_l904_l923_l917_DUPLICATE_74fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l920_l904_l923_l917_DUPLICATE_74fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l920_l904_l923_l917_DUPLICATE_74fb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l920_l904_l923_l917_DUPLICATE_74fb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l904_c2_d47e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l904_c2_d47e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l904_c2_d47e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l904_c2_d47e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l925_c30_66df_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l923_c7_0425] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_cond;
     result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_return_output := result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- n8_MUX[uxn_opcodes_h_l923_c7_0425] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l923_c7_0425_cond <= VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_cond;
     n8_MUX_uxn_opcodes_h_l923_c7_0425_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_iftrue;
     n8_MUX_uxn_opcodes_h_l923_c7_0425_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_return_output := n8_MUX_uxn_opcodes_h_l923_c7_0425_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l923_c7_0425] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l923_c7_0425] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l923_c7_0425] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_return_output;

     -- t8_MUX[uxn_opcodes_h_l920_c7_94ca] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l920_c7_94ca_cond <= VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_cond;
     t8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue;
     t8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output := t8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l923_c7_0425] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse := VAR_n8_MUX_uxn_opcodes_h_l923_c7_0425_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l923_c7_0425_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l923_c7_0425_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l923_c7_0425_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l923_c7_0425_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l923_c7_0425_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;
     -- t8_MUX[uxn_opcodes_h_l917_c7_722f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l917_c7_722f_cond <= VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_cond;
     t8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue;
     t8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_return_output := t8_MUX_uxn_opcodes_h_l917_c7_722f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l920_c7_94ca] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;

     -- n8_MUX[uxn_opcodes_h_l920_c7_94ca] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l920_c7_94ca_cond <= VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_cond;
     n8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue;
     n8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output := n8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l920_c7_94ca] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_cond;
     result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_return_output := result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l920_c7_94ca] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l920_c7_94ca] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l920_c7_94ca] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l920_c7_94ca_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l917_c7_722f_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l917_c7_722f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_return_output;

     -- t8_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     t8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     t8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := t8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- n8_MUX[uxn_opcodes_h_l917_c7_722f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l917_c7_722f_cond <= VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_cond;
     n8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_iftrue;
     n8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_return_output := n8_MUX_uxn_opcodes_h_l917_c7_722f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l917_c7_722f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l917_c7_722f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l917_c7_722f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_return_output := result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l917_c7_722f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l917_c7_722f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l917_c7_722f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l917_c7_722f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l917_c7_722f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l917_c7_722f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l917_c7_722f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- n8_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     n8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     n8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := n8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l904_c2_d47e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l904_c2_d47e_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l932_l900_DUPLICATE_eb2d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l932_l900_DUPLICATE_eb2d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l904_c2_d47e_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l904_c2_d47e_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l932_l900_DUPLICATE_eb2d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l932_l900_DUPLICATE_eb2d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
