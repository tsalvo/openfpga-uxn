-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sth2_0CLK_55b6500a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth2_0CLK_55b6500a;
architecture arch of sth2_0CLK_55b6500a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2436_c6_7d5e]
signal BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2436_c2_16f6]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2449_c11_8c95]
signal BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2449_c7_6c22]
signal t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2449_c7_6c22]
signal t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2449_c7_6c22]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2449_c7_6c22]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2449_c7_6c22]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2449_c7_6c22]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2449_c7_6c22]
signal result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2449_c7_6c22]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2452_c11_eab9]
signal BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2452_c7_c7a8]
signal t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(7 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2452_c7_c7a8]
signal t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2452_c7_c7a8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2452_c7_c7a8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2452_c7_c7a8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2452_c7_c7a8]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2452_c7_c7a8]
signal result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2452_c7_c7a8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2454_c30_2111]
signal sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2456_c11_ba2c]
signal BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2456_c7_c9fc]
signal t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2456_c7_c9fc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2456_c7_c9fc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2456_c7_c9fc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2456_c7_c9fc]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2456_c7_c9fc]
signal result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2456_c7_c9fc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2464_c11_7bd5]
signal BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2464_c7_3052]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2464_c7_3052]
signal result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2464_c7_3052]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2464_c7_3052]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_188e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_ram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e
BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_left,
BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_right,
BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6
t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6
t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6
result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6
result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6
result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6
result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95
BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_left,
BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_right,
BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22
t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_cond,
t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue,
t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse,
t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22
t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_cond,
t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue,
t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse,
t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22
result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22
result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22
result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_cond,
result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22
result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9
BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_left,
BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_right,
BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8
t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond,
t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue,
t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse,
t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8
t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond,
t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue,
t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse,
t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8
result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8
result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8
result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2454_c30_2111
sp_relative_shift_uxn_opcodes_h_l2454_c30_2111 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_ins,
sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_x,
sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_y,
sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c
BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_left,
BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_right,
BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc
t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond,
t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue,
t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse,
t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc
result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc
result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc
result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc
result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5
BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_left,
BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_right,
BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052
result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052
result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_cond,
result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052
result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output,
 t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output,
 t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output,
 t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output,
 t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output,
 t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output,
 sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output,
 t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2441_c3_cae4 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2446_c3_6ddd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2450_c3_0474 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2461_c3_2d0a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2459_c3_9d6d : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2465_c3_2db0 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2466_c3_4e38 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2452_l2436_l2449_l2464_DUPLICATE_af3d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_e6cf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2449_l2464_DUPLICATE_f4a0_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_8ff1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2452_l2456_l2449_l2464_DUPLICATE_4c39_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2452_l2464_DUPLICATE_85ea_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2432_l2471_DUPLICATE_a817_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2459_c3_9d6d := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2459_c3_9d6d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2461_c3_2d0a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2461_c3_2d0a;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2441_c3_cae4 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2441_c3_cae4;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2450_c3_0474 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2450_c3_0474;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2446_c3_6ddd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2446_c3_6ddd;
     VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2465_c3_2db0 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2465_c3_2db0;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2466_c3_4e38 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2466_c3_4e38;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_left := VAR_phase;
     VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse := t16_low;
     -- sp_relative_shift[uxn_opcodes_h_l2454_c30_2111] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_ins;
     sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_x;
     sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_return_output := sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2452_l2464_DUPLICATE_85ea LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2452_l2464_DUPLICATE_85ea_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2452_c11_eab9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2449_c11_8c95] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_left;
     BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output := BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2449_l2464_DUPLICATE_f4a0 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2449_l2464_DUPLICATE_f4a0_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2452_l2436_l2449_l2464_DUPLICATE_af3d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2452_l2436_l2449_l2464_DUPLICATE_af3d_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2456_c11_ba2c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_e6cf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_e6cf_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2464_c11_7bd5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2436_c6_7d5e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_8ff1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_8ff1_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2452_l2456_l2449_l2464_DUPLICATE_4c39 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2452_l2456_l2449_l2464_DUPLICATE_4c39_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2436_c6_7d5e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2449_c11_8c95_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2452_c11_eab9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2456_c11_ba2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2464_c11_7bd5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2449_l2464_DUPLICATE_f4a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2449_l2464_DUPLICATE_f4a0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2452_l2456_l2449_l2464_DUPLICATE_4c39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2452_l2456_l2449_l2464_DUPLICATE_4c39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2452_l2456_l2449_l2464_DUPLICATE_4c39_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2452_l2456_l2449_l2464_DUPLICATE_4c39_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_8ff1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_8ff1_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_8ff1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_e6cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_e6cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2452_l2456_l2449_DUPLICATE_e6cf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2452_l2464_DUPLICATE_85ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2452_l2464_DUPLICATE_85ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2452_l2436_l2449_l2464_DUPLICATE_af3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2452_l2436_l2449_l2464_DUPLICATE_af3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2452_l2436_l2449_l2464_DUPLICATE_af3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2452_l2436_l2449_l2464_DUPLICATE_af3d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2436_c2_16f6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2454_c30_2111_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2452_c7_c7a8] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond;
     t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output := t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2464_c7_3052] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2464_c7_3052] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2464_c7_3052] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_return_output := result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2456_c7_c9fc] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2456_c7_c9fc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2456_c7_c9fc] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond;
     t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output := t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2464_c7_3052] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2464_c7_3052_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2464_c7_3052_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2464_c7_3052_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2464_c7_3052_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2456_c7_c9fc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2452_c7_c7a8] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2456_c7_c9fc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2452_c7_c7a8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2449_c7_6c22] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_cond;
     t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output := t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2452_c7_c7a8] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond;
     t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output := t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2456_c7_c9fc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2456_c7_c9fc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2456_c7_c9fc_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;
     -- t16_low_MUX[uxn_opcodes_h_l2449_c7_6c22] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_cond;
     t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output := t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2452_c7_c7a8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2449_c7_6c22] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2452_c7_c7a8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2452_c7_c7a8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2449_c7_6c22] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2452_c7_c7a8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2452_c7_c7a8_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2449_c7_6c22] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2449_c7_6c22] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output := result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2449_c7_6c22] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2449_c7_6c22] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2449_c7_6c22_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2436_c2_16f6] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output := result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2432_l2471_DUPLICATE_a817 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2432_l2471_DUPLICATE_a817_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_188e(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2436_c2_16f6_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2432_l2471_DUPLICATE_a817_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2432_l2471_DUPLICATE_a817_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
