-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity div_0CLK_09f6f009 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end div_0CLK_09f6f009;
architecture arch of div_0CLK_09f6f009 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2078_c6_d554]
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal t8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal n8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2078_c2_58a0]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2091_c11_f397]
signal BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2091_c7_f103]
signal t8_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2091_c7_f103]
signal n8_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2091_c7_f103]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2091_c7_f103]
signal result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2091_c7_f103]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2091_c7_f103]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2091_c7_f103]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2094_c11_52ae]
signal BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2094_c7_6de9]
signal t8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2094_c7_6de9]
signal n8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2094_c7_6de9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2094_c7_6de9]
signal result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2094_c7_6de9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2094_c7_6de9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2094_c7_6de9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2097_c11_997a]
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2097_c7_1f63]
signal n8_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2097_c7_1f63]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2097_c7_1f63]
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2097_c7_1f63]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2097_c7_1f63]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2097_c7_1f63]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2099_c30_b623]
signal sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2102_c21_299b]
signal BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_return_output : unsigned(0 downto 0);

-- BIN_OP_DIV[uxn_opcodes_h_l2102_c35_e6df]
signal BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_left : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_right : unsigned(7 downto 0);
signal BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_return_output : unsigned(7 downto 0);

-- MUX[uxn_opcodes_h_l2102_c21_5173]
signal MUX_uxn_opcodes_h_l2102_c21_5173_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2102_c21_5173_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2102_c21_5173_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2102_c21_5173_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554
BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_left,
BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_right,
BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output);

-- t8_MUX_uxn_opcodes_h_l2078_c2_58a0
t8_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
t8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- n8_MUX_uxn_opcodes_h_l2078_c2_58a0
n8_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
n8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0
result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0
result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0
result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397
BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_left,
BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_right,
BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output);

-- t8_MUX_uxn_opcodes_h_l2091_c7_f103
t8_MUX_uxn_opcodes_h_l2091_c7_f103 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2091_c7_f103_cond,
t8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue,
t8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse,
t8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output);

-- n8_MUX_uxn_opcodes_h_l2091_c7_f103
n8_MUX_uxn_opcodes_h_l2091_c7_f103 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2091_c7_f103_cond,
n8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue,
n8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse,
n8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103
result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103
result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_cond,
result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103
result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103
result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae
BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_left,
BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_right,
BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output);

-- t8_MUX_uxn_opcodes_h_l2094_c7_6de9
t8_MUX_uxn_opcodes_h_l2094_c7_6de9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond,
t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue,
t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse,
t8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output);

-- n8_MUX_uxn_opcodes_h_l2094_c7_6de9
n8_MUX_uxn_opcodes_h_l2094_c7_6de9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond,
n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue,
n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse,
n8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9
result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9
result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a
BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_left,
BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_right,
BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output);

-- n8_MUX_uxn_opcodes_h_l2097_c7_1f63
n8_MUX_uxn_opcodes_h_l2097_c7_1f63 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2097_c7_1f63_cond,
n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue,
n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse,
n8_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_cond,
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2099_c30_b623
sp_relative_shift_uxn_opcodes_h_l2099_c30_b623 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_ins,
sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_x,
sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_y,
sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b
BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_left,
BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_right,
BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_return_output);

-- BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df
BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df : entity work.BIN_OP_DIV_uint8_t_uint8_t_0CLK_a148083c port map (
BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_left,
BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_right,
BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_return_output);

-- MUX_uxn_opcodes_h_l2102_c21_5173
MUX_uxn_opcodes_h_l2102_c21_5173 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2102_c21_5173_cond,
MUX_uxn_opcodes_h_l2102_c21_5173_iftrue,
MUX_uxn_opcodes_h_l2102_c21_5173_iffalse,
MUX_uxn_opcodes_h_l2102_c21_5173_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output,
 t8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 n8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output,
 t8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output,
 n8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output,
 t8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output,
 n8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output,
 n8_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output,
 sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_return_output,
 BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_return_output,
 MUX_uxn_opcodes_h_l2102_c21_5173_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2083_c3_3943 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2088_c3_33bb : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2092_c3_700a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2101_c3_2ffa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2102_c21_5173_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2102_c21_5173_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2102_c21_5173_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_return_output : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2102_c21_5173_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2091_l2094_l2078_l2097_DUPLICATE_f450_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_a0ac_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_ccf3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_0ff8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2094_l2097_DUPLICATE_8603_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2074_l2106_DUPLICATE_6bcd_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2101_c3_2ffa := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2101_c3_2ffa;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2092_c3_700a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2092_c3_700a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2088_c3_33bb := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2088_c3_33bb;
     VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_y := resize(to_signed(-1, 2), 4);
     VAR_MUX_uxn_opcodes_h_l2102_c21_5173_iftrue := resize(to_unsigned(0, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_right := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2083_c3_3943 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2083_c3_3943;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_left := VAR_phase;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_right := t8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_left := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse := t8;
     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2091_c11_f397] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_left;
     BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output := BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2078_c6_d554] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_left;
     BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output := BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2102_c21_299b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_a0ac LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_a0ac_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_ccf3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_ccf3_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2097_c11_997a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2094_l2097_DUPLICATE_8603 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2094_l2097_DUPLICATE_8603_return_output := result.stack_address_sp_offset;

     -- BIN_OP_DIV[uxn_opcodes_h_l2102_c35_e6df] LATENCY=0
     -- Inputs
     BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_left <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_left;
     BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_right <= VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_right;
     -- Outputs
     VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_return_output := BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2091_l2094_l2078_l2097_DUPLICATE_f450 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2091_l2094_l2078_l2097_DUPLICATE_f450_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2094_c11_52ae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_left;
     BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output := BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l2099_c30_b623] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_ins;
     sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_x;
     sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_return_output := sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_0ff8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_0ff8_return_output := result.is_stack_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_MUX_uxn_opcodes_h_l2102_c21_5173_iffalse := VAR_BIN_OP_DIV_uxn_opcodes_h_l2102_c35_e6df_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c6_d554_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2091_c11_f397_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_52ae_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2097_c11_997a_return_output;
     VAR_MUX_uxn_opcodes_h_l2102_c21_5173_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2102_c21_299b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_ccf3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_ccf3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_ccf3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_a0ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_a0ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_a0ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_0ff8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_0ff8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2091_l2094_l2097_DUPLICATE_0ff8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2094_l2097_DUPLICATE_8603_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2094_l2097_DUPLICATE_8603_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2091_l2094_l2078_l2097_DUPLICATE_f450_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2091_l2094_l2078_l2097_DUPLICATE_f450_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2091_l2094_l2078_l2097_DUPLICATE_f450_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2091_l2094_l2078_l2097_DUPLICATE_f450_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2078_c2_58a0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2099_c30_b623_return_output;
     -- result_is_vram_write_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- n8_MUX[uxn_opcodes_h_l2097_c7_1f63] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2097_c7_1f63_cond <= VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_cond;
     n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue;
     n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output := n8_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2097_c7_1f63] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2097_c7_1f63] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2097_c7_1f63] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2097_c7_1f63] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- MUX[uxn_opcodes_h_l2102_c21_5173] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2102_c21_5173_cond <= VAR_MUX_uxn_opcodes_h_l2102_c21_5173_cond;
     MUX_uxn_opcodes_h_l2102_c21_5173_iftrue <= VAR_MUX_uxn_opcodes_h_l2102_c21_5173_iftrue;
     MUX_uxn_opcodes_h_l2102_c21_5173_iffalse <= VAR_MUX_uxn_opcodes_h_l2102_c21_5173_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2102_c21_5173_return_output := MUX_uxn_opcodes_h_l2102_c21_5173_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2094_c7_6de9] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond <= VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond;
     t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue;
     t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output := t8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue := VAR_MUX_uxn_opcodes_h_l2102_c21_5173_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2097_c7_1f63] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output := result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2094_c7_6de9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2094_c7_6de9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;

     -- t8_MUX[uxn_opcodes_h_l2091_c7_f103] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2091_c7_f103_cond <= VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_cond;
     t8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue;
     t8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output := t8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2094_c7_6de9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2094_c7_6de9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_cond;
     n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue;
     n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output := n8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2094_c7_6de9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2097_c7_1f63_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;
     -- n8_MUX[uxn_opcodes_h_l2091_c7_f103] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2091_c7_f103_cond <= VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_cond;
     n8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue;
     n8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output := n8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;

     -- t8_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := t8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2091_c7_f103] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2091_c7_f103] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2091_c7_f103] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2094_c7_6de9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2091_c7_f103] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2094_c7_6de9_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;
     -- n8_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := n8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2091_c7_f103] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_return_output := result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2091_c7_f103_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2078_c2_58a0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2074_l2106_DUPLICATE_6bcd LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2074_l2106_DUPLICATE_6bcd_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2078_c2_58a0_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2074_l2106_DUPLICATE_6bcd_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l2074_l2106_DUPLICATE_6bcd_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
