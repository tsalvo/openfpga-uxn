-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_16;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out uint8_t_array_16_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_return_output : unsigned(0 downto 0);

-- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce]
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_cond : unsigned(0 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iftrue : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iffalse : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_return_output : unsigned(0 downto 0);

-- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1]
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_cond : unsigned(0 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iftrue : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iffalse : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_return_output : unsigned(0 downto 0);

-- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8]
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_cond : unsigned(0 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iftrue : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iffalse : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_return_output : unsigned(0 downto 0);

-- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e]
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_cond : unsigned(0 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iftrue : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iffalse : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_return_output : unsigned(0 downto 0);

-- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94]
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_cond : unsigned(0 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iftrue : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iffalse : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_return_output : unsigned(0 downto 0);

-- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79]
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_cond : unsigned(0 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iftrue : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iffalse : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_return_output : unsigned(0 downto 0);

-- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11]
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_cond : unsigned(0 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iftrue : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iffalse : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_return_output : unsigned(0 downto 0);

-- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29]
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_cond : unsigned(0 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iftrue : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iffalse : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_afcb( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_array_16_t is
 
  variable base : uint8_t_array_16_t; 
  variable return_output : uint8_t_array_16_t;
begin
      base.data(2) := ref_toks_0;
      base.data(8) := ref_toks_1;
      base.data(5) := ref_toks_2;
      base.data(11) := ref_toks_3;
      base.data(14) := ref_toks_4;
      base.data(3) := ref_toks_5;
      base.data(0) := ref_toks_6;
      base.data(6) := ref_toks_7;
      base.data(9) := ref_toks_8;
      base.data(15) := ref_toks_9;
      base.data(12) := ref_toks_10;
      base.data(1) := ref_toks_11;
      base.data(4) := ref_toks_12;
      base.data(10) := ref_toks_13;
      base.data(7) := ref_toks_14;
      base.data(13) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_return_output);

-- rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_cond,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iftrue,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iffalse,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_return_output);

-- rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_cond,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iftrue,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iffalse,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_return_output);

-- rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_cond,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iftrue,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iffalse,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_return_output);

-- rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_cond,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iftrue,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iffalse,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_return_output);

-- rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_cond,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iftrue,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iffalse,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_return_output);

-- rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_cond,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iftrue,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iffalse,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_return_output);

-- rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_cond,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iftrue,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iffalse,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_return_output);

-- rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_cond,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iftrue,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iffalse,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_return_output,
 rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_return_output,
 rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_return_output,
 rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_return_output,
 rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_return_output,
 rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_return_output,
 rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_return_output,
 rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_return_output,
 rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_16;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : uint8_t_array_16_t;
 variable VAR_base : uint8_t_16;
 variable VAR_rv : uint8_t_array_16_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_c27e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_7963_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_a056_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_2084_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_c71b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_d6c2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_7a80_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_1c30_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_8754_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_6c2a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_24fa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_fb02_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_d956_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c16_9309_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c15_cc4e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_ff52_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_afcb_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_5ae3_return_output : uint8_t_array_16_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_right := to_unsigned(14, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_right := to_unsigned(12, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_right := to_unsigned(13, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_right := to_unsigned(15, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_right := to_unsigned(11, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_right := to_unsigned(10, 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iftrue := VAR_elem_val;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iftrue := VAR_elem_val;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iftrue := VAR_elem_val;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iftrue := VAR_elem_val;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iftrue := VAR_elem_val;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iftrue := VAR_elem_val;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iftrue := VAR_elem_val;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iftrue := VAR_elem_val;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_left := VAR_var_dim_0;
     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_11_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_2084] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_2084_return_output := VAR_ref_toks_0(11);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_fb02] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_fb02_return_output := VAR_ref_toks_0(1);

     -- CONST_REF_RD_uint8_t_uint8_t_16_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_a056] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_a056_return_output := VAR_ref_toks_0(5);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_9_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_8754] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_8754_return_output := VAR_ref_toks_0(9);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_c27e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_c27e_return_output := VAR_ref_toks_0(2);

     -- CONST_REF_RD_uint8_t_uint8_t_16_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c15_cc4e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c15_cc4e_return_output := VAR_ref_toks_0(7);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_15_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_6c2a] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_6c2a_return_output := VAR_ref_toks_0(15);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_10_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c16_9309] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c16_9309_return_output := VAR_ref_toks_0(10);

     -- CONST_REF_RD_uint8_t_uint8_t_16_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_d6c2] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_d6c2_return_output := VAR_ref_toks_0(3);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_1c30] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_1c30_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_16_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_7a80] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_7a80_return_output := VAR_ref_toks_0(0);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_13_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_ff52] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_ff52_return_output := VAR_ref_toks_0(13);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_d956] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_d956_return_output := VAR_ref_toks_0(4);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_8_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_7963] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_7963_return_output := VAR_ref_toks_0(8);

     -- CONST_REF_RD_uint8_t_uint8_t_16_12_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_24fa] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_24fa_return_output := VAR_ref_toks_0(12);

     -- CONST_REF_RD_uint8_t_uint8_t_16_14_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_c71b] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_c71b_return_output := VAR_ref_toks_0(14);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_return_output;

     -- Submodule level 1
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_c691_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_b131_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_caad_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_4de7_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_fb7c_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_fffe_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_9899_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_16de_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_3018_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_3d03_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_4a2c_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_122d_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_eef3_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_c551_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_48e7_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_97aa_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_7a80_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c16_9309_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_2084_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_24fa_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_ff52_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c16_c71b_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c16_6c2a_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c15_fb02_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c15_c27e_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c15_d6c2_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_d956_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_a056_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_1c30_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c15_cc4e_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_7963_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_8754_return_output;
     -- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29] LATENCY=0
     -- Inputs
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_cond <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_cond;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iftrue;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_iffalse;
     -- Outputs
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_return_output := rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_return_output;

     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_return_output;

     -- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce] LATENCY=0
     -- Inputs
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_cond <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_cond;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iftrue;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_iffalse;
     -- Outputs
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_return_output := rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_return_output;

     -- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94] LATENCY=0
     -- Inputs
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_cond <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_cond;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iftrue;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_iffalse;
     -- Outputs
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_return_output := rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_return_output;

     -- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8] LATENCY=0
     -- Inputs
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_cond <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_cond;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iftrue;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_iffalse;
     -- Outputs
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_return_output := rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_return_output;

     -- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e] LATENCY=0
     -- Inputs
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_cond <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_cond;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iftrue;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_iffalse;
     -- Outputs
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_return_output := rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_return_output;

     -- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11] LATENCY=0
     -- Inputs
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_cond <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_cond;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iftrue;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_iffalse;
     -- Outputs
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_return_output := rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_return_output;

     -- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79] LATENCY=0
     -- Inputs
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_cond <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_cond;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iftrue;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_iffalse;
     -- Outputs
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_return_output := rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_return_output;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_return_output;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_return_output;

     -- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1] LATENCY=0
     -- Inputs
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_cond <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_cond;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iftrue;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_iffalse;
     -- Outputs
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_return_output := rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_afcb[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_5ae3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_afcb_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_5ae3_return_output := CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_afcb(
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_8b22_return_output,
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_42ce_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_914e_return_output,
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_76f1_return_output,
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_76e8_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_adfb_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_588f_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_56c5_return_output,
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_015e_return_output,
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_fc94_return_output,
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_7f79_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_73e4_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_25b4_return_output,
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_9e11_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_ca25_return_output,
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_4f29_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_afcb_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_5ae3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
