-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity ovr_0CLK_61914e8d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_61914e8d;
architecture arch of ovr_0CLK_61914e8d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l297_c6_f605]
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l297_c2_1eec]
signal n8_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l297_c2_1eec]
signal t8_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_1eec]
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l310_c11_932e]
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l310_c7_2c1b]
signal n8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l310_c7_2c1b]
signal t8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_2c1b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l310_c7_2c1b]
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_2c1b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_2c1b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_2c1b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l313_c11_6c2c]
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l313_c7_2bfd]
signal n8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l313_c7_2bfd]
signal t8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_2bfd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l313_c7_2bfd]
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_2bfd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_2bfd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_2bfd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l315_c30_5044]
signal sp_relative_shift_uxn_opcodes_h_l315_c30_5044_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_5044_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_5044_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l315_c30_5044_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l320_c11_6521]
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l320_c7_e087]
signal n8_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l320_c7_e087_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_e087]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_e087]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_e087]
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l320_c7_e087]
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l326_c11_5643]
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_dfcd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_dfcd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l326_c7_dfcd]
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_ee25( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605
BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_left,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_right,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output);

-- n8_MUX_uxn_opcodes_h_l297_c2_1eec
n8_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
n8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
n8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
n8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- t8_MUX_uxn_opcodes_h_l297_c2_1eec
t8_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
t8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
t8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
t8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec
result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e
BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_left,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_right,
BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output);

-- n8_MUX_uxn_opcodes_h_l310_c7_2c1b
n8_MUX_uxn_opcodes_h_l310_c7_2c1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond,
n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue,
n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse,
n8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output);

-- t8_MUX_uxn_opcodes_h_l310_c7_2c1b
t8_MUX_uxn_opcodes_h_l310_c7_2c1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond,
t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue,
t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse,
t8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b
result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_cond,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c
BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_left,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_right,
BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output);

-- n8_MUX_uxn_opcodes_h_l313_c7_2bfd
n8_MUX_uxn_opcodes_h_l313_c7_2bfd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond,
n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue,
n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse,
n8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output);

-- t8_MUX_uxn_opcodes_h_l313_c7_2bfd
t8_MUX_uxn_opcodes_h_l313_c7_2bfd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond,
t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue,
t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse,
t8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd
result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_cond,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output);

-- sp_relative_shift_uxn_opcodes_h_l315_c30_5044
sp_relative_shift_uxn_opcodes_h_l315_c30_5044 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l315_c30_5044_ins,
sp_relative_shift_uxn_opcodes_h_l315_c30_5044_x,
sp_relative_shift_uxn_opcodes_h_l315_c30_5044_y,
sp_relative_shift_uxn_opcodes_h_l315_c30_5044_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521
BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_left,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_right,
BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output);

-- n8_MUX_uxn_opcodes_h_l320_c7_e087
n8_MUX_uxn_opcodes_h_l320_c7_e087 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l320_c7_e087_cond,
n8_MUX_uxn_opcodes_h_l320_c7_e087_iftrue,
n8_MUX_uxn_opcodes_h_l320_c7_e087_iffalse,
n8_MUX_uxn_opcodes_h_l320_c7_e087_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087
result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_cond,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643
BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_left,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_right,
BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd
result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_cond,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output,
 n8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 t8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output,
 n8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output,
 t8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output,
 n8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output,
 t8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output,
 sp_relative_shift_uxn_opcodes_h_l315_c30_5044_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output,
 n8_MUX_uxn_opcodes_h_l320_c7_e087_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_8983 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_e167 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_31bd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_7113 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l321_c3_ca12 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_26d4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_dd2e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_dfcd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_41d7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_ccd1_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_8c4a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l320_l310_l326_l313_DUPLICATE_5f63_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l332_l293_DUPLICATE_5ff5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_right := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_8983 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l302_c3_8983;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_31bd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l311_c3_31bd;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_7113 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l317_c3_7113;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_e167 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l307_c3_e167;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l321_c3_ca12 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l321_c3_ca12;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_dd2e := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l327_c3_dd2e;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_26d4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l323_c3_26d4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l320_c11_6521] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_left;
     BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output := BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_1eec_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l326_c11_5643] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_left;
     BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output := BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_41d7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_41d7_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_1eec_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_1eec_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l310_c11_932e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_left;
     BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output := BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l297_c6_f605] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_left;
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output := BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_ccd1 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_ccd1_return_output := result.sp_relative_shift;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l326_c7_dfcd] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_dfcd_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l313_c11_6c2c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_left;
     BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output := BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_1eec_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l320_l310_l326_l313_DUPLICATE_5f63 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l320_l310_l326_l313_DUPLICATE_5f63_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_8c4a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_8c4a_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l315_c30_5044] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l315_c30_5044_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_ins;
     sp_relative_shift_uxn_opcodes_h_l315_c30_5044_x <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_x;
     sp_relative_shift_uxn_opcodes_h_l315_c30_5044_y <= VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_return_output := sp_relative_shift_uxn_opcodes_h_l315_c30_5044_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_f605_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l310_c11_932e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l313_c11_6c2c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l320_c11_6521_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l326_c11_5643_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_ccd1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l320_l310_DUPLICATE_ccd1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l320_l310_l326_l313_DUPLICATE_5f63_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l320_l310_l326_l313_DUPLICATE_5f63_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l320_l310_l326_l313_DUPLICATE_5f63_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l320_l310_l326_l313_DUPLICATE_5f63_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_8c4a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l310_l313_DUPLICATE_8c4a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_41d7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_41d7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l310_l326_DUPLICATE_41d7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l297_c2_1eec_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l297_c2_1eec_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l297_c2_1eec_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l297_c2_1eec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l326_c7_dfcd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l315_c30_5044_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l326_c7_dfcd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output := result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l326_c7_dfcd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output;

     -- t8_MUX[uxn_opcodes_h_l313_c7_2bfd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond;
     t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue;
     t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output := t8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l320_c7_e087] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l313_c7_2bfd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- n8_MUX[uxn_opcodes_h_l320_c7_e087] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l320_c7_e087_cond <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_cond;
     n8_MUX_uxn_opcodes_h_l320_c7_e087_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_iftrue;
     n8_MUX_uxn_opcodes_h_l320_c7_e087_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_return_output := n8_MUX_uxn_opcodes_h_l320_c7_e087_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l326_c7_dfcd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l320_c7_e087_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l320_c7_e087_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l326_c7_dfcd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l320_c7_e087] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_cond;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_return_output := result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l313_c7_2bfd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;

     -- n8_MUX[uxn_opcodes_h_l313_c7_2bfd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_cond;
     n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue;
     n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output := n8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;

     -- t8_MUX[uxn_opcodes_h_l310_c7_2c1b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond;
     t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue;
     t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output := t8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l320_c7_e087] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l310_c7_2c1b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l320_c7_e087] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l320_c7_e087_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l320_c7_e087_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l320_c7_e087_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_t8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l310_c7_2c1b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;

     -- n8_MUX[uxn_opcodes_h_l310_c7_2c1b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_cond;
     n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue;
     n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output := n8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;

     -- t8_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     t8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     t8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := t8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l313_c7_2bfd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l313_c7_2bfd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output := result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l313_c7_2bfd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_n8_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l313_c7_2bfd_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l310_c7_2c1b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;

     -- n8_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     n8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     n8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := n8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l310_c7_2c1b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output := result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l310_c7_2c1b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l310_c7_2c1b_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_1eec] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l332_l293_DUPLICATE_5ff5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l332_l293_DUPLICATE_5ff5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_ee25(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l297_c2_1eec_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l297_c2_1eec_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l332_l293_DUPLICATE_5ff5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_ee25_uxn_opcodes_h_l332_l293_DUPLICATE_5ff5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
