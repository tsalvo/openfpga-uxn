-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 41
entity jmp2_0CLK_0b1ee796 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jmp2_0CLK_0b1ee796;
architecture arch of jmp2_0CLK_0b1ee796 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l606_c6_5a14]
signal BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l606_c1_aca3]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l606_c2_74cb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l606_c2_74cb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l606_c2_74cb]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l606_c2_74cb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l606_c2_74cb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l606_c2_74cb]
signal result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l606_c2_74cb]
signal t16_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l607_c3_0457[uxn_opcodes_h_l607_c3_0457]
signal printf_uxn_opcodes_h_l607_c3_0457_uxn_opcodes_h_l607_c3_0457_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l611_c11_8ec7]
signal BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l611_c7_30a1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l611_c7_30a1]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l611_c7_30a1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l611_c7_30a1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l611_c7_30a1]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l611_c7_30a1]
signal result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l611_c7_30a1]
signal t16_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l614_c11_f183]
signal BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l614_c7_62ec]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l614_c7_62ec]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l614_c7_62ec]
signal result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l614_c7_62ec]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l614_c7_62ec]
signal result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l614_c7_62ec]
signal t16_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l616_c3_d681]
signal CONST_SL_8_uxn_opcodes_h_l616_c3_d681_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l616_c3_d681_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l618_c11_078c]
signal BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l618_c7_e867]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l618_c7_e867]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l618_c7_e867]
signal result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l618_c7_e867]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l618_c7_e867]
signal result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(15 downto 0);

-- t16_MUX[uxn_opcodes_h_l618_c7_e867]
signal t16_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l619_c3_b2ce]
signal BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l621_c30_81a3]
signal sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l625_c11_fb23]
signal BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l625_c7_24ea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l625_c7_24ea]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l625_c7_24ea]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_4c49( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : signed;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.sp_relative_shift := ref_toks_2;
      base.is_pc_updated := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_sp_shift := ref_toks_5;
      base.u16_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14
BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_left,
BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_right,
BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb
result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb
result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb
result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb
result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb
result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_cond,
result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_return_output);

-- t16_MUX_uxn_opcodes_h_l606_c2_74cb
t16_MUX_uxn_opcodes_h_l606_c2_74cb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l606_c2_74cb_cond,
t16_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue,
t16_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse,
t16_MUX_uxn_opcodes_h_l606_c2_74cb_return_output);

-- printf_uxn_opcodes_h_l607_c3_0457_uxn_opcodes_h_l607_c3_0457
printf_uxn_opcodes_h_l607_c3_0457_uxn_opcodes_h_l607_c3_0457 : entity work.printf_uxn_opcodes_h_l607_c3_0457_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l607_c3_0457_uxn_opcodes_h_l607_c3_0457_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7
BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_left,
BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_right,
BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1
result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1
result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1
result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1
result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1
result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_cond,
result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_return_output);

-- t16_MUX_uxn_opcodes_h_l611_c7_30a1
t16_MUX_uxn_opcodes_h_l611_c7_30a1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l611_c7_30a1_cond,
t16_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue,
t16_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse,
t16_MUX_uxn_opcodes_h_l611_c7_30a1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183
BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_left,
BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_right,
BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec
result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec
result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec
result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec
result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec
result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_cond,
result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_return_output);

-- t16_MUX_uxn_opcodes_h_l614_c7_62ec
t16_MUX_uxn_opcodes_h_l614_c7_62ec : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l614_c7_62ec_cond,
t16_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue,
t16_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse,
t16_MUX_uxn_opcodes_h_l614_c7_62ec_return_output);

-- CONST_SL_8_uxn_opcodes_h_l616_c3_d681
CONST_SL_8_uxn_opcodes_h_l616_c3_d681 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l616_c3_d681_x,
CONST_SL_8_uxn_opcodes_h_l616_c3_d681_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c
BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_left,
BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_right,
BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867
result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867
result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867
result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867
result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867
result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_cond,
result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_return_output);

-- t16_MUX_uxn_opcodes_h_l618_c7_e867
t16_MUX_uxn_opcodes_h_l618_c7_e867 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l618_c7_e867_cond,
t16_MUX_uxn_opcodes_h_l618_c7_e867_iftrue,
t16_MUX_uxn_opcodes_h_l618_c7_e867_iffalse,
t16_MUX_uxn_opcodes_h_l618_c7_e867_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce
BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_left,
BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_right,
BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_return_output);

-- sp_relative_shift_uxn_opcodes_h_l621_c30_81a3
sp_relative_shift_uxn_opcodes_h_l621_c30_81a3 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_ins,
sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_x,
sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_y,
sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23
BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_left,
BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_right,
BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea
result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea
result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea
result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
 t16_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_return_output,
 t16_MUX_uxn_opcodes_h_l611_c7_30a1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_return_output,
 t16_MUX_uxn_opcodes_h_l614_c7_62ec_return_output,
 CONST_SL_8_uxn_opcodes_h_l616_c3_d681_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_return_output,
 t16_MUX_uxn_opcodes_h_l618_c7_e867_return_output,
 BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_return_output,
 sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l608_c3_6aea : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l607_c3_0457_uxn_opcodes_h_l607_c3_0457_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l612_c3_7ca2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l611_c7_30a1_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l616_c3_d681_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l616_c3_d681_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_e12b_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_6ace_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_9fbb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_a354_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l614_l618_l611_l625_DUPLICATE_9145_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l619_l615_DUPLICATE_bbf9_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4c49_uxn_opcodes_h_l631_l602_DUPLICATE_3576_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_y := resize(to_signed(-2, 3), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l608_c3_6aea := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l608_c3_6aea;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue := to_unsigned(1, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l612_c3_7ca2 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l612_c3_7ca2;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_iffalse := t16;
     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_a354 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_a354_return_output := result.u16_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_e12b LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_e12b_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l618_c11_078c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_left;
     BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output := BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_6ace LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_6ace_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l614_c11_f183] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_left;
     BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output := BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l611_c11_8ec7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_left;
     BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output := BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_9fbb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_9fbb_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l621_c30_81a3] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_ins;
     sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_x <= VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_x;
     sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_y <= VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_return_output := sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l611_c7_30a1] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l611_c7_30a1_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l606_c6_5a14] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_left;
     BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output := BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l614_l618_l611_l625_DUPLICATE_9145 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l614_l618_l611_l625_DUPLICATE_9145_return_output := result.is_opc_done;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l619_l615_DUPLICATE_bbf9 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l619_l615_DUPLICATE_bbf9_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l625_c11_fb23] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_left;
     BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output := BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l606_c6_5a14_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l611_c11_8ec7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l614_c11_f183_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l618_c11_078c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l625_c11_fb23_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l619_l615_DUPLICATE_bbf9_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l616_c3_d681_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l619_l615_DUPLICATE_bbf9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_e12b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_e12b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_e12b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_e12b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_a354_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_a354_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_a354_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l614_l606_l618_l611_DUPLICATE_a354_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l614_l618_l611_l625_DUPLICATE_9145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l614_l618_l611_l625_DUPLICATE_9145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l614_l618_l611_l625_DUPLICATE_9145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l614_l618_l611_l625_DUPLICATE_9145_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_6ace_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_6ace_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_6ace_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_6ace_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_9fbb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_9fbb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_9fbb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l614_l606_l611_l625_DUPLICATE_9fbb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l611_c7_30a1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l621_c30_81a3_return_output;
     -- CONST_SL_8[uxn_opcodes_h_l616_c3_d681] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l616_c3_d681_x <= VAR_CONST_SL_8_uxn_opcodes_h_l616_c3_d681_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l616_c3_d681_return_output := CONST_SL_8_uxn_opcodes_h_l616_c3_d681_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l625_c7_24ea] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l619_c3_b2ce] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_left;
     BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_return_output := BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l618_c7_e867] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l606_c1_aca3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l625_c7_24ea] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l611_c7_30a1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l625_c7_24ea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l619_c3_b2ce_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l616_c3_d681_return_output;
     VAR_printf_uxn_opcodes_h_l607_c3_0457_uxn_opcodes_h_l607_c3_0457_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l606_c1_aca3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l625_c7_24ea_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l625_c7_24ea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l625_c7_24ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l618_c7_e867] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l618_c7_e867] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l618_c7_e867] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l618_c7_e867] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_cond;
     result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_return_output := result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_return_output;

     -- printf_uxn_opcodes_h_l607_c3_0457[uxn_opcodes_h_l607_c3_0457] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l607_c3_0457_uxn_opcodes_h_l607_c3_0457_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l607_c3_0457_uxn_opcodes_h_l607_c3_0457_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t16_MUX[uxn_opcodes_h_l618_c7_e867] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l618_c7_e867_cond <= VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_cond;
     t16_MUX_uxn_opcodes_h_l618_c7_e867_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_iftrue;
     t16_MUX_uxn_opcodes_h_l618_c7_e867_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_return_output := t16_MUX_uxn_opcodes_h_l618_c7_e867_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l606_c2_74cb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l614_c7_62ec] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l618_c7_e867_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l618_c7_e867_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l618_c7_e867_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l618_c7_e867_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse := VAR_t16_MUX_uxn_opcodes_h_l618_c7_e867_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l614_c7_62ec] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;

     -- t16_MUX[uxn_opcodes_h_l614_c7_62ec] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l614_c7_62ec_cond <= VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_cond;
     t16_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue;
     t16_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_return_output := t16_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l614_c7_62ec] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_cond;
     result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_return_output := result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l614_c7_62ec] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l614_c7_62ec] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l611_c7_30a1] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse := VAR_t16_MUX_uxn_opcodes_h_l614_c7_62ec_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l606_c2_74cb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l611_c7_30a1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l611_c7_30a1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l611_c7_30a1] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_cond;
     result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_return_output := result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l611_c7_30a1] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;

     -- t16_MUX[uxn_opcodes_h_l611_c7_30a1] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l611_c7_30a1_cond <= VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_cond;
     t16_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_iftrue;
     t16_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_return_output := t16_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse := VAR_t16_MUX_uxn_opcodes_h_l611_c7_30a1_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l606_c2_74cb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output;

     -- t16_MUX[uxn_opcodes_h_l606_c2_74cb] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l606_c2_74cb_cond <= VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_cond;
     t16_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue;
     t16_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_return_output := t16_MUX_uxn_opcodes_h_l606_c2_74cb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l606_c2_74cb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l606_c2_74cb] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_cond;
     result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_return_output := result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l606_c2_74cb] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_return_output;

     -- Submodule level 6
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l606_c2_74cb_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4c49_uxn_opcodes_h_l631_l602_DUPLICATE_3576 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4c49_uxn_opcodes_h_l631_l602_DUPLICATE_3576_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4c49(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l606_c2_74cb_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l606_c2_74cb_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4c49_uxn_opcodes_h_l631_l602_DUPLICATE_3576_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4c49_uxn_opcodes_h_l631_l602_DUPLICATE_3576_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
