-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 55
entity lit_0CLK_3220bbf1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lit_0CLK_3220bbf1;
architecture arch of lit_0CLK_3220bbf1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l206_c6_8cba]
signal BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l206_c1_7675]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(7 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(15 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : signed(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);

-- result_is_ram_read_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l206_c2_e22a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l206_c2_e22a]
signal tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l207_c3_5531[uxn_opcodes_h_l207_c3_5531]
signal printf_uxn_opcodes_h_l207_c3_5531_uxn_opcodes_h_l207_c3_5531_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l212_c11_a65a]
signal BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(7 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(15 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_pc_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);

-- result_is_ram_read_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l212_c7_2667]
signal result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l212_c7_2667]
signal tmp8_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l217_c11_333a]
signal BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l217_c7_42b1]
signal result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(7 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l217_c7_42b1]
signal result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(15 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l217_c7_42b1]
signal result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l217_c7_42b1]
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l217_c7_42b1]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(7 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l217_c7_42b1]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(0 downto 0);

-- result_is_ram_read_MUX[uxn_opcodes_h_l217_c7_42b1]
signal result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l217_c7_42b1]
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l217_c7_42b1]
signal tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l220_c11_52f0]
signal BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output : unsigned(0 downto 0);

-- result_is_ram_read_MUX[uxn_opcodes_h_l220_c7_2877]
signal result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(0 downto 0);
signal result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l220_c7_2877]
signal result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(7 downto 0);

-- result_pc_MUX[uxn_opcodes_h_l220_c7_2877]
signal result_pc_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(15 downto 0);
signal result_pc_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(15 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l220_c7_2877]
signal result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l220_c7_2877]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l220_c7_2877]
signal result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l220_c7_2877]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l220_c7_2877]
signal tmp8_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(7 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l224_c15_e091]
signal BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_left : unsigned(15 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_return_output : unsigned(16 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l226_c11_154a]
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output : unsigned(0 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l226_c7_dd89]
signal result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l226_c7_dd89]
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l226_c7_dd89]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l226_c7_dd89]
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l226_c7_dd89]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l232_c11_218e]
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l232_c7_9be7]
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l232_c7_9be7]
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_2e50( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_value := ref_toks_1;
      base.ram_addr := ref_toks_2;
      base.pc := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_sp_shift := ref_toks_8;
      base.is_ram_read := ref_toks_9;
      base.is_opc_done := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba
BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_left,
BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_right,
BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a
result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_pc_MUX_uxn_opcodes_h_l206_c2_e22a
result_pc_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- tmp8_MUX_uxn_opcodes_h_l206_c2_e22a
tmp8_MUX_uxn_opcodes_h_l206_c2_e22a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_cond,
tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue,
tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse,
tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

-- printf_uxn_opcodes_h_l207_c3_5531_uxn_opcodes_h_l207_c3_5531
printf_uxn_opcodes_h_l207_c3_5531_uxn_opcodes_h_l207_c3_5531 : entity work.printf_uxn_opcodes_h_l207_c3_5531_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l207_c3_5531_uxn_opcodes_h_l207_c3_5531_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a
BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_left,
BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_right,
BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667
result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- result_pc_MUX_uxn_opcodes_h_l212_c7_2667
result_pc_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_pc_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- tmp8_MUX_uxn_opcodes_h_l212_c7_2667
tmp8_MUX_uxn_opcodes_h_l212_c7_2667 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l212_c7_2667_cond,
tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iftrue,
tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iffalse,
tmp8_MUX_uxn_opcodes_h_l212_c7_2667_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a
BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_left,
BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_right,
BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1
result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- result_pc_MUX_uxn_opcodes_h_l217_c7_42b1
result_pc_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- tmp8_MUX_uxn_opcodes_h_l217_c7_42b1
tmp8_MUX_uxn_opcodes_h_l217_c7_42b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_cond,
tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue,
tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse,
tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0
BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_left,
BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_right,
BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output);

-- result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_cond,
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iftrue,
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iffalse,
result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877
result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_cond,
result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_return_output);

-- result_pc_MUX_uxn_opcodes_h_l220_c7_2877
result_pc_MUX_uxn_opcodes_h_l220_c7_2877 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_pc_MUX_uxn_opcodes_h_l220_c7_2877_cond,
result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iftrue,
result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iffalse,
result_pc_MUX_uxn_opcodes_h_l220_c7_2877_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_return_output);

-- tmp8_MUX_uxn_opcodes_h_l220_c7_2877
tmp8_MUX_uxn_opcodes_h_l220_c7_2877 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l220_c7_2877_cond,
tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iftrue,
tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iffalse,
tmp8_MUX_uxn_opcodes_h_l220_c7_2877_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091
BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091 : entity work.BIN_OP_PLUS_uint16_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_left,
BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_right,
BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a
BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_left,
BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_right,
BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89
result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_cond,
result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e
BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_left,
BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_right,
BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 previous_ram_read,
 -- Registers
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 result_pc_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 tmp8_MUX_uxn_opcodes_h_l212_c7_2667_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output,
 result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_return_output,
 result_pc_MUX_uxn_opcodes_h_l220_c7_2877_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_return_output,
 tmp8_MUX_uxn_opcodes_h_l220_c7_2877_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l209_c3_6277 : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l206_c2_e22a_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l207_c3_5531_uxn_opcodes_h_l207_c3_5531_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l212_c7_2667_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(15 downto 0);
 variable VAR_result_pc_uxn_opcodes_h_l224_c3_ff2c : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(15 downto 0);
 variable VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_return_output : unsigned(16 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l229_c3_1935 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_a11f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_d14d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l220_l212_l206_l217_DUPLICATE_0088_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l212_l217_l232_l206_DUPLICATE_17e5_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_e893_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l226_l212_l206_l217_DUPLICATE_2e45_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l220_l206_l217_DUPLICATE_3d04_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l226_l212_l217_l232_DUPLICATE_3c6d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2e50_uxn_opcodes_h_l201_l237_DUPLICATE_7ff1_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_right := to_unsigned(3, 2);
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_right := to_unsigned(4, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l229_c3_1935 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l229_c3_1935;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l209_c3_6277 := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l209_c3_6277;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iftrue := VAR_CLOCK_ENABLE;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_left := VAR_pc;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := VAR_pc;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_left := VAR_phase;
     VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iftrue := VAR_previous_ram_read;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iffalse := tmp8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l212_l217_l232_l206_DUPLICATE_17e5 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l212_l217_l232_l206_DUPLICATE_17e5_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_e893 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_e893_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l220_l206_l217_DUPLICATE_3d04 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l220_l206_l217_DUPLICATE_3d04_return_output := result.is_ram_read;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_a11f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_a11f_return_output := result.stack_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l220_c11_52f0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_left;
     BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output := BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l206_c6_8cba] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_left;
     BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output := BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l226_c11_154a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_left;
     BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output := BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output;

     -- result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l212_c7_2667_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l226_l212_l217_l232_DUPLICATE_3c6d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l226_l212_l217_l232_DUPLICATE_3c6d_return_output := result.is_opc_done;

     -- BIN_OP_PLUS[uxn_opcodes_h_l224_c15_e091] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_left;
     BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_return_output := BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_return_output;

     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l206_c2_e22a_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l220_l212_l206_l217_DUPLICATE_0088 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l220_l212_l206_l217_DUPLICATE_0088_return_output := result.pc;

     -- BIN_OP_EQ[uxn_opcodes_h_l232_c11_218e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_left;
     BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_return_output := BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l217_c11_333a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_left;
     BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output := BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l212_c11_a65a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_left;
     BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output := BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l226_l212_l206_l217_DUPLICATE_2e45 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l226_l212_l206_l217_DUPLICATE_2e45_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_d14d LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_d14d_return_output := result.ram_addr;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l206_c6_8cba_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l212_c11_a65a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l217_c11_333a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l220_c11_52f0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l226_c11_154a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l232_c11_218e_return_output;
     VAR_result_pc_uxn_opcodes_h_l224_c3_ff2c := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l224_c15_e091_return_output, 16);
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l220_l212_l206_l217_DUPLICATE_0088_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l220_l212_l206_l217_DUPLICATE_0088_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l220_l212_l206_l217_DUPLICATE_0088_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_pc_d41d_uxn_opcodes_h_l220_l212_l206_l217_DUPLICATE_0088_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_d14d_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l206_l217_DUPLICATE_d14d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l226_l212_l217_l232_DUPLICATE_3c6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l226_l212_l217_l232_DUPLICATE_3c6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l226_l212_l217_l232_DUPLICATE_3c6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l226_l212_l217_l232_DUPLICATE_3c6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l220_l226_l212_l217_l232_DUPLICATE_3c6d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l226_l212_l206_l217_DUPLICATE_2e45_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l226_l212_l206_l217_DUPLICATE_2e45_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l226_l212_l206_l217_DUPLICATE_2e45_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l226_l212_l206_l217_DUPLICATE_2e45_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l220_l206_l217_DUPLICATE_3d04_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l220_l206_l217_DUPLICATE_3d04_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_read_d41d_uxn_opcodes_h_l220_l206_l217_DUPLICATE_3d04_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l212_l217_l232_l206_DUPLICATE_17e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l212_l217_l232_l206_DUPLICATE_17e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l212_l217_l232_l206_DUPLICATE_17e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l212_l217_l232_l206_DUPLICATE_17e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l220_l212_l217_l232_l206_DUPLICATE_17e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_e893_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_e893_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_e893_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_e893_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_e893_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_a11f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_a11f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_a11f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_a11f_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l220_l226_l212_l217_l206_DUPLICATE_a11f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_is_sp_shift_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l212_c7_2667_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l206_c2_e22a_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iftrue := VAR_result_pc_uxn_opcodes_h_l224_c3_ff2c;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l226_c7_dd89] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_cond;
     result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_return_output := result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- result_is_ram_read_MUX[uxn_opcodes_h_l220_c7_2877] LATENCY=0
     -- Inputs
     result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_cond <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_cond;
     result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iftrue <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iftrue;
     result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iffalse <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_iffalse;
     -- Outputs
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_return_output := result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l226_c7_dd89] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l220_c7_2877] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l220_c7_2877_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_cond;
     result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iftrue;
     result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_return_output := result_pc_MUX_uxn_opcodes_h_l220_c7_2877_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l226_c7_dd89] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l232_c7_9be7] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l220_c7_2877] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l220_c7_2877_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_cond;
     tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iftrue;
     tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_return_output := tmp8_MUX_uxn_opcodes_h_l220_c7_2877_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l232_c7_9be7] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l206_c1_7675] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l207_c3_5531_uxn_opcodes_h_l207_c3_5531_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l206_c1_7675_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l232_c7_9be7_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_result_is_ram_read_MUX_uxn_opcodes_h_l220_c7_2877_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l232_c7_9be7_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l220_c7_2877_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l220_c7_2877_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l226_c7_dd89] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l220_c7_2877] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_cond;
     result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_return_output := result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l220_c7_2877] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l220_c7_2877] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_return_output;

     -- result_is_ram_read_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- printf_uxn_opcodes_h_l207_c3_5531[uxn_opcodes_h_l207_c3_5531] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l207_c3_5531_uxn_opcodes_h_l207_c3_5531_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l207_c3_5531_uxn_opcodes_h_l207_c3_5531_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- tmp8_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l226_c7_dd89] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l220_c7_2877_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_is_ram_read_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l226_c7_dd89_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l220_c7_2877_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l220_c7_2877_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l220_c7_2877] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_pc_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- result_is_ram_read_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_return_output := tmp8_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l220_c7_2877] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l220_c7_2877_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_is_ram_read_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l220_c7_2877_return_output;
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_pc_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     -- result_is_ram_read_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_pc_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l217_c7_42b1] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l217_c7_42b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l212_c7_2667] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l212_c7_2667_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l206_c2_e22a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_2e50_uxn_opcodes_h_l201_l237_DUPLICATE_7ff1 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2e50_uxn_opcodes_h_l201_l237_DUPLICATE_7ff1_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_2e50(
     result,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_pc_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_is_ram_read_MUX_uxn_opcodes_h_l206_c2_e22a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l206_c2_e22a_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2e50_uxn_opcodes_h_l201_l237_DUPLICATE_7ff1_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_2e50_uxn_opcodes_h_l201_l237_DUPLICATE_7ff1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
