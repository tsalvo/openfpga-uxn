-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 41
entity ovr_0CLK_282a76ca is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ovr_0CLK_282a76ca;
architecture arch of ovr_0CLK_282a76ca is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l297_c6_4dad]
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l297_c2_5a3c]
signal n8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l297_c2_5a3c]
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_5a3c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_5a3c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_5a3c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_5a3c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l297_c2_5a3c]
signal t8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l304_c11_aa2e]
signal BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l304_c7_5ad0]
signal n8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l304_c7_5ad0]
signal result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l304_c7_5ad0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l304_c7_5ad0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l304_c7_5ad0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l304_c7_5ad0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l304_c7_5ad0]
signal t8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l307_c11_5bfc]
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l307_c7_d467]
signal n8_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l307_c7_d467]
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_d467]
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_d467]
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_d467]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l307_c7_d467]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l307_c7_d467]
signal t8_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l310_c30_18b8]
signal sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l315_c11_8b55]
signal BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l315_c7_1a06]
signal n8_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l315_c7_1a06]
signal result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l315_c7_1a06]
signal result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l315_c7_1a06]
signal result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l315_c7_1a06]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l315_c7_1a06]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l321_c11_beb2]
signal BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l321_c7_38e9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l321_c7_38e9]
signal result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l321_c7_38e9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l321_c7_38e9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l325_c11_624b]
signal BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l325_c7_b71c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l325_c7_b71c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad
BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_left,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_right,
BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output);

-- n8_MUX_uxn_opcodes_h_l297_c2_5a3c
n8_MUX_uxn_opcodes_h_l297_c2_5a3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond,
n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue,
n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse,
n8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c
result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_cond,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output);

-- t8_MUX_uxn_opcodes_h_l297_c2_5a3c
t8_MUX_uxn_opcodes_h_l297_c2_5a3c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond,
t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue,
t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse,
t8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e
BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_left,
BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_right,
BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output);

-- n8_MUX_uxn_opcodes_h_l304_c7_5ad0
n8_MUX_uxn_opcodes_h_l304_c7_5ad0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond,
n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue,
n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse,
n8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0
result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_cond,
result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0
result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0
result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0
result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output);

-- t8_MUX_uxn_opcodes_h_l304_c7_5ad0
t8_MUX_uxn_opcodes_h_l304_c7_5ad0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond,
t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue,
t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse,
t8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc
BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_left,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_right,
BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output);

-- n8_MUX_uxn_opcodes_h_l307_c7_d467
n8_MUX_uxn_opcodes_h_l307_c7_d467 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l307_c7_d467_cond,
n8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue,
n8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse,
n8_MUX_uxn_opcodes_h_l307_c7_d467_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467
result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_cond,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467
result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_return_output);

-- t8_MUX_uxn_opcodes_h_l307_c7_d467
t8_MUX_uxn_opcodes_h_l307_c7_d467 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l307_c7_d467_cond,
t8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue,
t8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse,
t8_MUX_uxn_opcodes_h_l307_c7_d467_return_output);

-- sp_relative_shift_uxn_opcodes_h_l310_c30_18b8
sp_relative_shift_uxn_opcodes_h_l310_c30_18b8 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_ins,
sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_x,
sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_y,
sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55
BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_left,
BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_right,
BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output);

-- n8_MUX_uxn_opcodes_h_l315_c7_1a06
n8_MUX_uxn_opcodes_h_l315_c7_1a06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l315_c7_1a06_cond,
n8_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue,
n8_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse,
n8_MUX_uxn_opcodes_h_l315_c7_1a06_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06
result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_cond,
result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2
BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_left,
BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_right,
BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9
result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9
result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_cond,
result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9
result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b
BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_left,
BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_right,
BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c
result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output,
 n8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
 t8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output,
 n8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output,
 t8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output,
 n8_MUX_uxn_opcodes_h_l307_c7_d467_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_return_output,
 t8_MUX_uxn_opcodes_h_l307_c7_d467_return_output,
 sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output,
 n8_MUX_uxn_opcodes_h_l315_c7_1a06_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l301_c3_5308 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_ac78 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l312_c3_bbc1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l318_c3_ae46 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l316_c3_3f95 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l322_c3_1a37 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l321_c7_38e9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l304_l321_DUPLICATE_a978_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l304_l297_l325_l321_l315_DUPLICATE_fbd6_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l297_l315_l304_DUPLICATE_3d81_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l304_l325_l321_l315_l307_DUPLICATE_a0cf_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l330_l293_DUPLICATE_1e04_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_ac78 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l305_c3_ac78;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l318_c3_ae46 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l318_c3_ae46;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l316_c3_3f95 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l316_c3_3f95;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l312_c3_bbc1 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l312_c3_bbc1;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l322_c3_1a37 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l322_c3_1a37;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l301_c3_5308 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l301_c3_5308;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse := n8;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l315_c11_8b55] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_left;
     BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output := BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l321_c7_38e9] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l321_c7_38e9_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l310_c30_18b8] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_ins;
     sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_x <= VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_x;
     sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_y <= VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_return_output := sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l304_l321_DUPLICATE_a978 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l304_l321_DUPLICATE_a978_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l297_l315_l304_DUPLICATE_3d81 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l297_l315_l304_DUPLICATE_3d81_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l297_c6_4dad] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_left;
     BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output := BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l307_c11_5bfc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_left;
     BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output := BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l304_l325_l321_l315_l307_DUPLICATE_a0cf LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l304_l325_l321_l315_l307_DUPLICATE_a0cf_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l325_c11_624b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_left;
     BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_return_output := BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l321_c11_beb2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_left;
     BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output := BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l304_l297_l325_l321_l315_DUPLICATE_fbd6 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l304_l297_l325_l321_l315_DUPLICATE_fbd6_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l304_c11_aa2e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_left;
     BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output := BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l297_c6_4dad_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l304_c11_aa2e_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l307_c11_5bfc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l315_c11_8b55_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l321_c11_beb2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l325_c11_624b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l297_l315_l304_DUPLICATE_3d81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l297_l315_l304_DUPLICATE_3d81_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l297_l315_l304_DUPLICATE_3d81_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l304_l325_l321_l315_l307_DUPLICATE_a0cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l304_l325_l321_l315_l307_DUPLICATE_a0cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l304_l325_l321_l315_l307_DUPLICATE_a0cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l304_l325_l321_l315_l307_DUPLICATE_a0cf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l304_l325_l321_l315_l307_DUPLICATE_a0cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l304_l297_l325_l321_l315_DUPLICATE_fbd6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l304_l297_l325_l321_l315_DUPLICATE_fbd6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l304_l297_l325_l321_l315_DUPLICATE_fbd6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l304_l297_l325_l321_l315_DUPLICATE_fbd6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l304_l297_l325_l321_l315_DUPLICATE_fbd6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l304_l321_DUPLICATE_a978_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l304_l321_DUPLICATE_a978_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l297_l304_l321_DUPLICATE_a978_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l321_c7_38e9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l310_c30_18b8_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l321_c7_38e9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_return_output;

     -- n8_MUX[uxn_opcodes_h_l315_c7_1a06] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l315_c7_1a06_cond <= VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_cond;
     n8_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue;
     n8_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_return_output := n8_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l315_c7_1a06] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l321_c7_38e9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_return_output := result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l325_c7_b71c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l325_c7_b71c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_return_output;

     -- t8_MUX[uxn_opcodes_h_l307_c7_d467] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l307_c7_d467_cond <= VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_cond;
     t8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue;
     t8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_return_output := t8_MUX_uxn_opcodes_h_l307_c7_d467_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse := VAR_n8_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l325_c7_b71c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l325_c7_b71c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l321_c7_38e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l321_c7_38e9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l307_c7_d467_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l315_c7_1a06] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_cond;
     result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_return_output := result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l321_c7_38e9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_return_output;

     -- n8_MUX[uxn_opcodes_h_l307_c7_d467] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l307_c7_d467_cond <= VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_cond;
     n8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_iftrue;
     n8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_return_output := n8_MUX_uxn_opcodes_h_l307_c7_d467_return_output;

     -- t8_MUX[uxn_opcodes_h_l304_c7_5ad0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond <= VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond;
     t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue;
     t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output := t8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l307_c7_d467] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l321_c7_38e9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l315_c7_1a06] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l307_c7_d467_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l321_c7_38e9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l321_c7_38e9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l307_c7_d467_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l304_c7_5ad0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l307_c7_d467] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_cond;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_return_output := result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l315_c7_1a06] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l315_c7_1a06] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;

     -- n8_MUX[uxn_opcodes_h_l304_c7_5ad0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond <= VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_cond;
     n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue;
     n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output := n8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;

     -- t8_MUX[uxn_opcodes_h_l297_c2_5a3c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond;
     t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue;
     t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output := t8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l307_c7_d467] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l315_c7_1a06_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l307_c7_d467_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l307_c7_d467_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l304_c7_5ad0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output := result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;

     -- n8_MUX[uxn_opcodes_h_l297_c2_5a3c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_cond;
     n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue;
     n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output := n8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l307_c7_d467] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l307_c7_d467] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l297_c2_5a3c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l304_c7_5ad0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l307_c7_d467_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l307_c7_d467_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l297_c2_5a3c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l304_c7_5ad0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l297_c2_5a3c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output := result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l304_c7_5ad0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l304_c7_5ad0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l297_c2_5a3c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l297_c2_5a3c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l330_l293_DUPLICATE_1e04 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l330_l293_DUPLICATE_1e04_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l297_c2_5a3c_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l330_l293_DUPLICATE_1e04_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l330_l293_DUPLICATE_1e04_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
