-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity eor_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end eor_0CLK_64d180f1;
architecture arch of eor_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1076_c6_62ed]
signal BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1076_c2_bbd3]
signal t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1089_c11_afb9]
signal BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1089_c7_a971]
signal n8_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1089_c7_a971]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1089_c7_a971]
signal result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1089_c7_a971]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1089_c7_a971]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1089_c7_a971]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1089_c7_a971]
signal t8_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1092_c11_56a6]
signal BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1092_c7_55bd]
signal n8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1092_c7_55bd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1092_c7_55bd]
signal result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1092_c7_55bd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1092_c7_55bd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1092_c7_55bd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1092_c7_55bd]
signal t8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1095_c11_ddca]
signal BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1095_c7_5878]
signal n8_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1095_c7_5878]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1095_c7_5878]
signal result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1095_c7_5878]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1095_c7_5878]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1095_c7_5878]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1097_c30_0c09]
signal sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_return_output : signed(3 downto 0);

-- BIN_OP_XOR[uxn_opcodes_h_l1100_c21_bd0a]
signal BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_left : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_right : unsigned(7 downto 0);
signal BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_vram_write := ref_toks_3;
      base.is_pc_updated := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.stack_address_sp_offset := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed
BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_left,
BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_right,
BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output);

-- n8_MUX_uxn_opcodes_h_l1076_c2_bbd3
n8_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- t8_MUX_uxn_opcodes_h_l1076_c2_bbd3
t8_MUX_uxn_opcodes_h_l1076_c2_bbd3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond,
t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue,
t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse,
t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9
BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_left,
BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_right,
BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output);

-- n8_MUX_uxn_opcodes_h_l1089_c7_a971
n8_MUX_uxn_opcodes_h_l1089_c7_a971 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1089_c7_a971_cond,
n8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue,
n8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse,
n8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971
result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971
result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_cond,
result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971
result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971
result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_return_output);

-- t8_MUX_uxn_opcodes_h_l1089_c7_a971
t8_MUX_uxn_opcodes_h_l1089_c7_a971 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1089_c7_a971_cond,
t8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue,
t8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse,
t8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6
BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_left,
BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_right,
BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output);

-- n8_MUX_uxn_opcodes_h_l1092_c7_55bd
n8_MUX_uxn_opcodes_h_l1092_c7_55bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond,
n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue,
n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse,
n8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd
result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd
result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_cond,
result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd
result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd
result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output);

-- t8_MUX_uxn_opcodes_h_l1092_c7_55bd
t8_MUX_uxn_opcodes_h_l1092_c7_55bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond,
t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue,
t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse,
t8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca
BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_left,
BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_right,
BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output);

-- n8_MUX_uxn_opcodes_h_l1095_c7_5878
n8_MUX_uxn_opcodes_h_l1095_c7_5878 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1095_c7_5878_cond,
n8_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue,
n8_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse,
n8_MUX_uxn_opcodes_h_l1095_c7_5878_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878
result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878
result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_cond,
result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878
result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878
result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09
sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_ins,
sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_x,
sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_y,
sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_return_output);

-- BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a
BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a : entity work.BIN_OP_XOR_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_left,
BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_right,
BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output,
 n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output,
 n8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_return_output,
 t8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output,
 n8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output,
 t8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output,
 n8_MUX_uxn_opcodes_h_l1095_c7_5878_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_return_output,
 sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_return_output,
 BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1081_c3_ad3e : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1086_c3_c849 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1090_c3_f428 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1099_c3_04c9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1089_l1092_l1076_l1095_DUPLICATE_1d45_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_e2ad_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_c8d5_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_11ac_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1092_l1095_DUPLICATE_7232_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1104_l1072_DUPLICATE_d05f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1081_c3_ad3e := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1081_c3_ad3e;
     VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_y := resize(to_signed(-1, 2), 4);
     VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1099_c3_04c9 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1099_c3_04c9;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1090_c3_f428 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1090_c3_f428;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1086_c3_c849 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1086_c3_c849;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_left := VAR_phase;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse := t8;
     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output := result.is_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1092_c11_56a6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1089_l1092_l1076_l1095_DUPLICATE_1d45 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1089_l1092_l1076_l1095_DUPLICATE_1d45_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_c8d5 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_c8d5_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1092_l1095_DUPLICATE_7232 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1092_l1095_DUPLICATE_7232_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1095_c11_ddca] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_left;
     BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output := BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output;

     -- BIN_OP_XOR[uxn_opcodes_h_l1100_c21_bd0a] LATENCY=0
     -- Inputs
     BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_left <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_left;
     BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_right <= VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_right;
     -- Outputs
     VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_return_output := BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_11ac LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_11ac_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_e2ad LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_e2ad_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l1097_c30_0c09] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_ins;
     sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_x;
     sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_return_output := sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1089_c11_afb9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1076_c6_62ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1076_c6_62ed_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1089_c11_afb9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1092_c11_56a6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1095_c11_ddca_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue := VAR_BIN_OP_XOR_uxn_opcodes_h_l1100_c21_bd0a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_c8d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_c8d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_c8d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_11ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_11ac_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_11ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_e2ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_e2ad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1089_l1092_l1095_DUPLICATE_e2ad_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1092_l1095_DUPLICATE_7232_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1092_l1095_DUPLICATE_7232_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1089_l1092_l1076_l1095_DUPLICATE_1d45_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1089_l1092_l1076_l1095_DUPLICATE_1d45_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1089_l1092_l1076_l1095_DUPLICATE_1d45_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1089_l1092_l1076_l1095_DUPLICATE_1d45_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1076_c2_bbd3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1097_c30_0c09_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1095_c7_5878] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1095_c7_5878] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1095_c7_5878_cond <= VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_cond;
     n8_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue;
     n8_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_return_output := n8_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1095_c7_5878] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1095_c7_5878] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_return_output := result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1095_c7_5878] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;

     -- t8_MUX[uxn_opcodes_h_l1092_c7_55bd] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond <= VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond;
     t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue;
     t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output := t8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1095_c7_5878] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1095_c7_5878_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;
     -- t8_MUX[uxn_opcodes_h_l1089_c7_a971] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1089_c7_a971_cond <= VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_cond;
     t8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue;
     t8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output := t8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;

     -- n8_MUX[uxn_opcodes_h_l1092_c7_55bd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond <= VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_cond;
     n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue;
     n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output := n8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1092_c7_55bd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1092_c7_55bd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1092_c7_55bd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1092_c7_55bd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1092_c7_55bd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output := result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1092_c7_55bd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1089_c7_a971] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_return_output := result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1089_c7_a971] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1089_c7_a971] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1089_c7_a971] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1089_c7_a971] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;

     -- t8_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1089_c7_a971] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1089_c7_a971_cond <= VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_cond;
     n8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_iftrue;
     n8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output := n8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1089_c7_a971_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;
     -- n8_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1076_c2_bbd3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1104_l1072_DUPLICATE_d05f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1104_l1072_DUPLICATE_d05f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1076_c2_bbd3_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1104_l1072_DUPLICATE_d05f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c5ea_uxn_opcodes_h_l1104_l1072_DUPLICATE_d05f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
