-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 37
entity dup_0CLK_6be78140 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end dup_0CLK_6be78140;
architecture arch of dup_0CLK_6be78140 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2616_c6_34c8]
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2616_c1_f12b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2616_c2_2d05]
signal t8_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2616_c2_2d05]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2616_c2_2d05]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2616_c2_2d05]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2616_c2_2d05]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2616_c2_2d05]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2616_c2_2d05]
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2617_c3_b0c6[uxn_opcodes_h_l2617_c3_b0c6]
signal printf_uxn_opcodes_h_l2617_c3_b0c6_uxn_opcodes_h_l2617_c3_b0c6_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2621_c11_0cc5]
signal BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2621_c7_7f10]
signal t8_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2621_c7_7f10]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2621_c7_7f10]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2621_c7_7f10]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2621_c7_7f10]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2621_c7_7f10]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2621_c7_7f10]
signal result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2624_c11_4e58]
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2624_c7_5391]
signal t8_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2624_c7_5391]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2624_c7_5391]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2624_c7_5391]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2624_c7_5391]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2624_c7_5391]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2624_c7_5391]
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2627_c30_169f]
signal sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2632_c11_e8f4]
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2632_c7_ab3a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2632_c7_ab3a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2632_c7_ab3a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2632_c7_ab3a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2632_c7_ab3a]
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2637_c11_4e44]
signal BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2637_c7_01dc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2637_c7_01dc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8
BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_left,
BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_right,
BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_return_output);

-- t8_MUX_uxn_opcodes_h_l2616_c2_2d05
t8_MUX_uxn_opcodes_h_l2616_c2_2d05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2616_c2_2d05_cond,
t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue,
t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse,
t8_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05
result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_cond,
result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output);

-- printf_uxn_opcodes_h_l2617_c3_b0c6_uxn_opcodes_h_l2617_c3_b0c6
printf_uxn_opcodes_h_l2617_c3_b0c6_uxn_opcodes_h_l2617_c3_b0c6 : entity work.printf_uxn_opcodes_h_l2617_c3_b0c6_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2617_c3_b0c6_uxn_opcodes_h_l2617_c3_b0c6_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5
BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_left,
BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_right,
BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output);

-- t8_MUX_uxn_opcodes_h_l2621_c7_7f10
t8_MUX_uxn_opcodes_h_l2621_c7_7f10 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2621_c7_7f10_cond,
t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue,
t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse,
t8_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10
result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10
result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10
result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10
result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10
result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_cond,
result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_left,
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_right,
BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output);

-- t8_MUX_uxn_opcodes_h_l2624_c7_5391
t8_MUX_uxn_opcodes_h_l2624_c7_5391 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2624_c7_5391_cond,
t8_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue,
t8_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse,
t8_MUX_uxn_opcodes_h_l2624_c7_5391_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_cond,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2627_c30_169f
sp_relative_shift_uxn_opcodes_h_l2627_c30_169f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_ins,
sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_x,
sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_y,
sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_left,
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_right,
BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44
BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_left,
BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_right,
BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_return_output,
 t8_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output,
 t8_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output,
 t8_MUX_uxn_opcodes_h_l2624_c7_5391_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_return_output,
 sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2618_c3_e0a0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2617_c3_b0c6_uxn_opcodes_h_l2617_c3_b0c6_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_f84d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2629_c3_b64e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2634_c3_acfd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2632_c7_ab3a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_89fd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2616_l2632_l2621_l2637_DUPLICATE_9827_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2624_l2616_l2621_DUPLICATE_0c64_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_0d7b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2632_l2621_l2637_DUPLICATE_5f34_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2642_l2612_DUPLICATE_17e9_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_y := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_f84d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2622_c3_f84d;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2634_c3_acfd := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2634_c3_acfd;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iffalse := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2629_c3_b64e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2629_c3_b64e;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2618_c3_e0a0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2618_c3_e0a0;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_right := to_unsigned(4, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l2627_c30_169f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_ins;
     sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_x;
     sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_return_output := sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_0d7b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_0d7b_return_output := result.u8_value;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2632_c7_ab3a] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2632_c7_ab3a_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2632_l2621_l2637_DUPLICATE_5f34 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2632_l2621_l2637_DUPLICATE_5f34_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2632_c11_e8f4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_left;
     BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output := BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2624_l2616_l2621_DUPLICATE_0c64 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2624_l2616_l2621_DUPLICATE_0c64_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_89fd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_89fd_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2637_c11_4e44] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_left;
     BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_return_output := BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2624_c11_4e58] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_left;
     BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output := BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2616_c6_34c8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2621_c11_0cc5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2616_l2632_l2621_l2637_DUPLICATE_9827 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2616_l2632_l2621_l2637_DUPLICATE_9827_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2616_c6_34c8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2621_c11_0cc5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2624_c11_4e58_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2632_c11_e8f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2637_c11_4e44_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2624_l2616_l2621_DUPLICATE_0c64_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2624_l2616_l2621_DUPLICATE_0c64_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2624_l2616_l2621_DUPLICATE_0c64_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2632_l2621_l2637_DUPLICATE_5f34_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2632_l2621_l2637_DUPLICATE_5f34_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2632_l2621_l2637_DUPLICATE_5f34_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2624_l2632_l2621_l2637_DUPLICATE_5f34_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_89fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_89fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_89fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2616_l2632_l2621_l2637_DUPLICATE_9827_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2616_l2632_l2621_l2637_DUPLICATE_9827_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2616_l2632_l2621_l2637_DUPLICATE_9827_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2616_l2632_l2621_l2637_DUPLICATE_9827_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_0d7b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_0d7b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2616_l2632_l2621_DUPLICATE_0d7b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2632_c7_ab3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2627_c30_169f_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2632_c7_ab3a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;

     -- t8_MUX[uxn_opcodes_h_l2624_c7_5391] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2624_c7_5391_cond <= VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_cond;
     t8_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue;
     t8_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_return_output := t8_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2632_c7_ab3a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2637_c7_01dc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2637_c7_01dc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2632_c7_ab3a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2616_c1_f12b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2624_c7_5391] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2617_c3_b0c6_uxn_opcodes_h_l2617_c3_b0c6_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2616_c1_f12b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2637_c7_01dc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2632_c7_ab3a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2624_c7_5391] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_return_output := result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2632_c7_ab3a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2624_c7_5391] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;

     -- printf_uxn_opcodes_h_l2617_c3_b0c6[uxn_opcodes_h_l2617_c3_b0c6] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2617_c3_b0c6_uxn_opcodes_h_l2617_c3_b0c6_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2617_c3_b0c6_uxn_opcodes_h_l2617_c3_b0c6_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2621_c7_7f10] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;

     -- t8_MUX[uxn_opcodes_h_l2621_c7_7f10] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2621_c7_7f10_cond <= VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_cond;
     t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue;
     t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output := t8_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2624_c7_5391] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2632_c7_ab3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2624_c7_5391] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2621_c7_7f10] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2616_c2_2d05] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2621_c7_7f10] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output := result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2624_c7_5391] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2621_c7_7f10] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;

     -- t8_MUX[uxn_opcodes_h_l2616_c2_2d05] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2616_c2_2d05_cond <= VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_cond;
     t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue;
     t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output := t8_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2624_c7_5391_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2616_c2_2d05] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2616_c2_2d05] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output := result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2621_c7_7f10] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2616_c2_2d05] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2621_c7_7f10] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2621_c7_7f10_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2616_c2_2d05] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2616_c2_2d05] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2642_l2612_DUPLICATE_17e9 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2642_l2612_DUPLICATE_17e9_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2616_c2_2d05_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2642_l2612_DUPLICATE_17e9_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2642_l2612_DUPLICATE_17e9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
