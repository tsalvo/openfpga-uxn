-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_46cced44 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_46cced44;
architecture arch of sft_0CLK_46cced44 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2213_c6_fdec]
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal n8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2213_c2_0c85]
signal t8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2226_c11_7376]
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2226_c7_9a41]
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2226_c7_9a41]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2226_c7_9a41]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2226_c7_9a41]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2226_c7_9a41]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2226_c7_9a41]
signal n8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2226_c7_9a41]
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2226_c7_9a41]
signal t8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2229_c11_2b3a]
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2229_c7_26ea]
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2229_c7_26ea]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2229_c7_26ea]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2229_c7_26ea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2229_c7_26ea]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2229_c7_26ea]
signal n8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2229_c7_26ea]
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2229_c7_26ea]
signal t8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2231_c30_eeaa]
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2233_c11_85ff]
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2233_c7_13d4]
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2233_c7_13d4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2233_c7_13d4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2233_c7_13d4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2233_c7_13d4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2233_c7_13d4]
signal n8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2233_c7_13d4]
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2236_c18_68d7]
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2236_c11_52e8]
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2236_c34_1c80]
signal CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2236_c11_98f2]
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_922a( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_pc_updated := ref_toks_6;
      base.is_opc_done := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_left,
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_right,
BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- n8_MUX_uxn_opcodes_h_l2213_c2_0c85
n8_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
n8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85
tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- t8_MUX_uxn_opcodes_h_l2213_c2_0c85
t8_MUX_uxn_opcodes_h_l2213_c2_0c85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond,
t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue,
t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse,
t8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_left,
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_right,
BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_cond,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output);

-- n8_MUX_uxn_opcodes_h_l2226_c7_9a41
n8_MUX_uxn_opcodes_h_l2226_c7_9a41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond,
n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue,
n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse,
n8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41
tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond,
tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue,
tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse,
tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output);

-- t8_MUX_uxn_opcodes_h_l2226_c7_9a41
t8_MUX_uxn_opcodes_h_l2226_c7_9a41 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond,
t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue,
t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse,
t8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_left,
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_right,
BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_cond,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output);

-- n8_MUX_uxn_opcodes_h_l2229_c7_26ea
n8_MUX_uxn_opcodes_h_l2229_c7_26ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond,
n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue,
n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse,
n8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea
tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond,
tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue,
tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse,
tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output);

-- t8_MUX_uxn_opcodes_h_l2229_c7_26ea
t8_MUX_uxn_opcodes_h_l2229_c7_26ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond,
t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue,
t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse,
t8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa
sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_ins,
sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_x,
sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_y,
sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_left,
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_right,
BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_cond,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output);

-- n8_MUX_uxn_opcodes_h_l2233_c7_13d4
n8_MUX_uxn_opcodes_h_l2233_c7_13d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond,
n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue,
n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse,
n8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4
tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond,
tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue,
tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse,
tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7
BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_left,
BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_right,
BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8
BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8 : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_left,
BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_right,
BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80
CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80 : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_x,
CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2
BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2 : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_left,
BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_right,
BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 n8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 t8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output,
 n8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output,
 tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output,
 t8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output,
 n8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output,
 tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output,
 t8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output,
 sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output,
 n8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output,
 tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_return_output,
 CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_921d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_9c1c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_8f15 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_e540 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_88c8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_c5ed_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_9aaf_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_7fca_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_410a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_6b90_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2209_l2243_DUPLICATE_29e5_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_right := to_unsigned(3, 2);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_921d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2223_c3_921d;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_y := resize(to_signed(-1, 2), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_88c8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2235_c3_88c8;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_8f15 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2227_c3_8f15;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_e540 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2238_c3_e540;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_right := to_unsigned(15, 8);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_9c1c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2218_c3_9c1c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_right := to_unsigned(2, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse := tmp8;
     -- BIN_OP_AND[uxn_opcodes_h_l2236_c18_68d7] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_left;
     BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_return_output := BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_9aaf LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_9aaf_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_410a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_410a_return_output := result.is_stack_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output := result.is_pc_updated;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l2231_c30_eeaa] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_ins;
     sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_x;
     sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_return_output := sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2233_c11_85ff] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_left;
     BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output := BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2229_c11_2b3a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2226_c11_7376] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_left;
     BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output := BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;

     -- CONST_SR_4[uxn_opcodes_h_l2236_c34_1c80] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_return_output := CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_6b90 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_6b90_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2213_c6_fdec] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_left;
     BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output := BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_c5ed LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_c5ed_return_output := result.u8_value;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_7fca LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_7fca_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2236_c18_68d7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2213_c6_fdec_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2226_c11_7376_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2229_c11_2b3a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2233_c11_85ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_9aaf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2233_l2226_DUPLICATE_9aaf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_7fca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_7fca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_7fca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_410a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_410a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2229_l2233_l2226_DUPLICATE_410a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_6b90_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2229_l2233_DUPLICATE_6b90_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_c5ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_c5ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_c5ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2229_l2213_l2233_l2226_DUPLICATE_c5ed_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_right := VAR_CONST_SR_4_uxn_opcodes_h_l2236_c34_1c80_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2213_c2_0c85_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2231_c30_eeaa_return_output;
     -- t8_MUX[uxn_opcodes_h_l2229_c7_26ea] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond;
     t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue;
     t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output := t8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;

     -- BIN_OP_SR[uxn_opcodes_h_l2236_c11_52e8] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_left;
     BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_return_output := BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- n8_MUX[uxn_opcodes_h_l2233_c7_13d4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond;
     n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue;
     n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output := n8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2233_c7_13d4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2233_c7_13d4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2233_c7_13d4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2233_c7_13d4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2236_c11_52e8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2229_c7_26ea] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2236_c11_98f2] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_left;
     BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_return_output := BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2229_c7_26ea] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2229_c7_26ea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;

     -- n8_MUX[uxn_opcodes_h_l2229_c7_26ea] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond;
     n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue;
     n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output := n8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2229_c7_26ea] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;

     -- t8_MUX[uxn_opcodes_h_l2226_c7_9a41] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond;
     t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue;
     t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output := t8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2236_c11_98f2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;
     -- t8_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := t8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2233_c7_13d4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output := result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2226_c7_9a41] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2226_c7_9a41] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2226_c7_9a41] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2226_c7_9a41] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2233_c7_13d4] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_cond;
     tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output := tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;

     -- n8_MUX[uxn_opcodes_h_l2226_c7_9a41] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond;
     n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue;
     n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output := n8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2233_c7_13d4_return_output;
     -- n8_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := n8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2229_c7_26ea] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output := result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2229_c7_26ea] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_cond;
     tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output := tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2229_c7_26ea_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2226_c7_9a41] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_cond;
     tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output := tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2226_c7_9a41] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output := result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2226_c7_9a41_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2213_c2_0c85] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_cond;
     tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output := tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2209_l2243_DUPLICATE_29e5 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2209_l2243_DUPLICATE_29e5_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_922a(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2213_c2_0c85_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2209_l2243_DUPLICATE_29e5_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_922a_uxn_opcodes_h_l2209_l2243_DUPLICATE_29e5_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
