-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 48
entity swp_0CLK_faaf4b1a is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp_0CLK_faaf4b1a;
architecture arch of swp_0CLK_faaf4b1a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2414_c6_0746]
signal BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2414_c1_42fd]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2414_c2_22af]
signal t8_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2414_c2_22af]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2414_c2_22af]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2414_c2_22af]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2414_c2_22af]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2414_c2_22af]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2414_c2_22af]
signal result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2414_c2_22af]
signal n8_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2415_c3_95d4[uxn_opcodes_h_l2415_c3_95d4]
signal printf_uxn_opcodes_h_l2415_c3_95d4_uxn_opcodes_h_l2415_c3_95d4_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2419_c11_e159]
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2419_c7_b91f]
signal t8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c7_b91f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2419_c7_b91f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c7_b91f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c7_b91f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c7_b91f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2419_c7_b91f]
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2419_c7_b91f]
signal n8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2422_c11_9380]
signal BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2422_c7_2d22]
signal t8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2422_c7_2d22]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2422_c7_2d22]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2422_c7_2d22]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2422_c7_2d22]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2422_c7_2d22]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2422_c7_2d22]
signal result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2422_c7_2d22]
signal n8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2425_c11_98af]
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c7_d17b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2425_c7_d17b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c7_d17b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c7_d17b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2425_c7_d17b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2425_c7_d17b]
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2425_c7_d17b]
signal n8_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2428_c30_b184]
signal sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2433_c11_a711]
signal BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2433_c7_ac88]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2433_c7_ac88]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2433_c7_ac88]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2433_c7_ac88]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2433_c7_ac88]
signal result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2438_c11_4104]
signal BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2438_c7_d360]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2438_c7_d360]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746
BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_left,
BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_right,
BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_return_output);

-- t8_MUX_uxn_opcodes_h_l2414_c2_22af
t8_MUX_uxn_opcodes_h_l2414_c2_22af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2414_c2_22af_cond,
t8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue,
t8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse,
t8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af
result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_cond,
result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

-- n8_MUX_uxn_opcodes_h_l2414_c2_22af
n8_MUX_uxn_opcodes_h_l2414_c2_22af : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2414_c2_22af_cond,
n8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue,
n8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse,
n8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

-- printf_uxn_opcodes_h_l2415_c3_95d4_uxn_opcodes_h_l2415_c3_95d4
printf_uxn_opcodes_h_l2415_c3_95d4_uxn_opcodes_h_l2415_c3_95d4 : entity work.printf_uxn_opcodes_h_l2415_c3_95d4_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2415_c3_95d4_uxn_opcodes_h_l2415_c3_95d4_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159
BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_left,
BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_right,
BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output);

-- t8_MUX_uxn_opcodes_h_l2419_c7_b91f
t8_MUX_uxn_opcodes_h_l2419_c7_b91f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond,
t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue,
t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse,
t8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f
result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output);

-- n8_MUX_uxn_opcodes_h_l2419_c7_b91f
n8_MUX_uxn_opcodes_h_l2419_c7_b91f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond,
n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue,
n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse,
n8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380
BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_left,
BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_right,
BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output);

-- t8_MUX_uxn_opcodes_h_l2422_c7_2d22
t8_MUX_uxn_opcodes_h_l2422_c7_2d22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond,
t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue,
t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse,
t8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22
result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_cond,
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output);

-- n8_MUX_uxn_opcodes_h_l2422_c7_2d22
n8_MUX_uxn_opcodes_h_l2422_c7_2d22 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond,
n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue,
n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse,
n8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_left,
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_right,
BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output);

-- n8_MUX_uxn_opcodes_h_l2425_c7_d17b
n8_MUX_uxn_opcodes_h_l2425_c7_d17b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2425_c7_d17b_cond,
n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue,
n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse,
n8_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2428_c30_b184
sp_relative_shift_uxn_opcodes_h_l2428_c30_b184 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_ins,
sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_x,
sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_y,
sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711
BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_left,
BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_right,
BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88
result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_cond,
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104
BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_left,
BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_right,
BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_return_output,
 t8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
 n8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output,
 t8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output,
 n8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output,
 t8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output,
 n8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output,
 n8_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output,
 sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2416_c3_1d97 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2415_c3_95d4_uxn_opcodes_h_l2415_c3_95d4_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2420_c3_c16c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_6f84 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2435_c3_9660 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_874c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2438_l2433_l2422_l2419_DUPLICATE_3d75_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2422_l2414_l2425_l2419_DUPLICATE_f21d_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_c2d2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2433_l2425_l2422_l2419_DUPLICATE_2663_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2433_DUPLICATE_2314_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2410_l2443_DUPLICATE_b8e3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_right := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2420_c3_c16c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2420_c3_c16c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_6f84 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2430_c3_6f84;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2416_c3_1d97 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2416_c3_1d97;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_right := to_unsigned(5, 3);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2435_c3_9660 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2435_c3_9660;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2438_l2433_l2422_l2419_DUPLICATE_3d75 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2438_l2433_l2422_l2419_DUPLICATE_3d75_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l2428_c30_b184] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_ins;
     sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_x;
     sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_return_output := sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2419_c11_e159] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_left;
     BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output := BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2425_c11_98af] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_left;
     BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output := BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2438_c11_4104] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_left;
     BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_return_output := BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2422_c11_9380] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_left;
     BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output := BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_c2d2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_c2d2_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2433_c11_a711] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_left;
     BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output := BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2433_l2425_l2422_l2419_DUPLICATE_2663 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2433_l2425_l2422_l2419_DUPLICATE_2663_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_874c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_874c_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2414_c6_0746] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_left;
     BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output := BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2433_DUPLICATE_2314 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2433_DUPLICATE_2314_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2422_l2414_l2425_l2419_DUPLICATE_f21d LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2422_l2414_l2425_l2419_DUPLICATE_f21d_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2414_c6_0746_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_e159_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2422_c11_9380_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2425_c11_98af_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2433_c11_a711_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2438_c11_4104_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2422_l2414_l2425_l2419_DUPLICATE_f21d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2422_l2414_l2425_l2419_DUPLICATE_f21d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2422_l2414_l2425_l2419_DUPLICATE_f21d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2422_l2414_l2425_l2419_DUPLICATE_f21d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2433_l2425_l2422_l2419_DUPLICATE_2663_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2433_l2425_l2422_l2419_DUPLICATE_2663_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2433_l2425_l2422_l2419_DUPLICATE_2663_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2433_l2425_l2422_l2419_DUPLICATE_2663_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2438_l2433_l2425_l2422_l2419_DUPLICATE_2663_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_874c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_874c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_874c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_874c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2438_l2433_l2422_l2419_DUPLICATE_3d75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2438_l2433_l2422_l2419_DUPLICATE_3d75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2438_l2433_l2422_l2419_DUPLICATE_3d75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2438_l2433_l2422_l2419_DUPLICATE_3d75_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2414_l2438_l2433_l2422_l2419_DUPLICATE_3d75_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2433_DUPLICATE_2314_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2422_l2433_DUPLICATE_2314_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_c2d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_c2d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_c2d2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2422_l2414_l2419_l2433_DUPLICATE_c2d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2428_c30_b184_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2438_c7_d360] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_return_output;

     -- t8_MUX[uxn_opcodes_h_l2422_c7_2d22] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond <= VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond;
     t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue;
     t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output := t8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;

     -- n8_MUX[uxn_opcodes_h_l2425_c7_d17b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2425_c7_d17b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_cond;
     n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue;
     n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output := n8_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2425_c7_d17b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2433_c7_ac88] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2433_c7_ac88] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output := result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2414_c1_42fd] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2433_c7_ac88] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2438_c7_d360] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2415_c3_95d4_uxn_opcodes_h_l2415_c3_95d4_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2414_c1_42fd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2438_c7_d360_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2438_c7_d360_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2425_c7_d17b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2419_c7_b91f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond;
     t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue;
     t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output := t8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2422_c7_2d22] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;

     -- n8_MUX[uxn_opcodes_h_l2422_c7_2d22] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond <= VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_cond;
     n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue;
     n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output := n8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;

     -- printf_uxn_opcodes_h_l2415_c3_95d4[uxn_opcodes_h_l2415_c3_95d4] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2415_c3_95d4_uxn_opcodes_h_l2415_c3_95d4_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2415_c3_95d4_uxn_opcodes_h_l2415_c3_95d4_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2425_c7_d17b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2425_c7_d17b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2433_c7_ac88] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2433_c7_ac88] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2433_c7_ac88_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2422_c7_2d22] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output := result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2425_c7_d17b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;

     -- n8_MUX[uxn_opcodes_h_l2419_c7_b91f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond <= VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_cond;
     n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue;
     n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output := n8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2414_c2_22af] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2414_c2_22af_cond <= VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_cond;
     t8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue;
     t8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output := t8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2425_c7_d17b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2422_c7_2d22] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c7_b91f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2422_c7_2d22] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2425_c7_d17b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c7_b91f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2422_c7_2d22] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2414_c2_22af] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2419_c7_b91f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2422_c7_2d22] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;

     -- n8_MUX[uxn_opcodes_h_l2414_c2_22af] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2414_c2_22af_cond <= VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_cond;
     n8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue;
     n8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output := n8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2419_c7_b91f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2422_c7_2d22_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2414_c2_22af] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_return_output := result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2414_c2_22af] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2414_c2_22af] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c7_b91f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c7_b91f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_b91f_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2414_c2_22af] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2414_c2_22af] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2410_l2443_DUPLICATE_b8e3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2410_l2443_DUPLICATE_b8e3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2414_c2_22af_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2414_c2_22af_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2410_l2443_DUPLICATE_b8e3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2410_l2443_DUPLICATE_b8e3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
