-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 134
entity uint8_mux128_0CLK_9347d63d is
port(
 sel : in unsigned(6 downto 0);
 in0 : in unsigned(7 downto 0);
 in1 : in unsigned(7 downto 0);
 in2 : in unsigned(7 downto 0);
 in3 : in unsigned(7 downto 0);
 in4 : in unsigned(7 downto 0);
 in5 : in unsigned(7 downto 0);
 in6 : in unsigned(7 downto 0);
 in7 : in unsigned(7 downto 0);
 in8 : in unsigned(7 downto 0);
 in9 : in unsigned(7 downto 0);
 in10 : in unsigned(7 downto 0);
 in11 : in unsigned(7 downto 0);
 in12 : in unsigned(7 downto 0);
 in13 : in unsigned(7 downto 0);
 in14 : in unsigned(7 downto 0);
 in15 : in unsigned(7 downto 0);
 in16 : in unsigned(7 downto 0);
 in17 : in unsigned(7 downto 0);
 in18 : in unsigned(7 downto 0);
 in19 : in unsigned(7 downto 0);
 in20 : in unsigned(7 downto 0);
 in21 : in unsigned(7 downto 0);
 in22 : in unsigned(7 downto 0);
 in23 : in unsigned(7 downto 0);
 in24 : in unsigned(7 downto 0);
 in25 : in unsigned(7 downto 0);
 in26 : in unsigned(7 downto 0);
 in27 : in unsigned(7 downto 0);
 in28 : in unsigned(7 downto 0);
 in29 : in unsigned(7 downto 0);
 in30 : in unsigned(7 downto 0);
 in31 : in unsigned(7 downto 0);
 in32 : in unsigned(7 downto 0);
 in33 : in unsigned(7 downto 0);
 in34 : in unsigned(7 downto 0);
 in35 : in unsigned(7 downto 0);
 in36 : in unsigned(7 downto 0);
 in37 : in unsigned(7 downto 0);
 in38 : in unsigned(7 downto 0);
 in39 : in unsigned(7 downto 0);
 in40 : in unsigned(7 downto 0);
 in41 : in unsigned(7 downto 0);
 in42 : in unsigned(7 downto 0);
 in43 : in unsigned(7 downto 0);
 in44 : in unsigned(7 downto 0);
 in45 : in unsigned(7 downto 0);
 in46 : in unsigned(7 downto 0);
 in47 : in unsigned(7 downto 0);
 in48 : in unsigned(7 downto 0);
 in49 : in unsigned(7 downto 0);
 in50 : in unsigned(7 downto 0);
 in51 : in unsigned(7 downto 0);
 in52 : in unsigned(7 downto 0);
 in53 : in unsigned(7 downto 0);
 in54 : in unsigned(7 downto 0);
 in55 : in unsigned(7 downto 0);
 in56 : in unsigned(7 downto 0);
 in57 : in unsigned(7 downto 0);
 in58 : in unsigned(7 downto 0);
 in59 : in unsigned(7 downto 0);
 in60 : in unsigned(7 downto 0);
 in61 : in unsigned(7 downto 0);
 in62 : in unsigned(7 downto 0);
 in63 : in unsigned(7 downto 0);
 in64 : in unsigned(7 downto 0);
 in65 : in unsigned(7 downto 0);
 in66 : in unsigned(7 downto 0);
 in67 : in unsigned(7 downto 0);
 in68 : in unsigned(7 downto 0);
 in69 : in unsigned(7 downto 0);
 in70 : in unsigned(7 downto 0);
 in71 : in unsigned(7 downto 0);
 in72 : in unsigned(7 downto 0);
 in73 : in unsigned(7 downto 0);
 in74 : in unsigned(7 downto 0);
 in75 : in unsigned(7 downto 0);
 in76 : in unsigned(7 downto 0);
 in77 : in unsigned(7 downto 0);
 in78 : in unsigned(7 downto 0);
 in79 : in unsigned(7 downto 0);
 in80 : in unsigned(7 downto 0);
 in81 : in unsigned(7 downto 0);
 in82 : in unsigned(7 downto 0);
 in83 : in unsigned(7 downto 0);
 in84 : in unsigned(7 downto 0);
 in85 : in unsigned(7 downto 0);
 in86 : in unsigned(7 downto 0);
 in87 : in unsigned(7 downto 0);
 in88 : in unsigned(7 downto 0);
 in89 : in unsigned(7 downto 0);
 in90 : in unsigned(7 downto 0);
 in91 : in unsigned(7 downto 0);
 in92 : in unsigned(7 downto 0);
 in93 : in unsigned(7 downto 0);
 in94 : in unsigned(7 downto 0);
 in95 : in unsigned(7 downto 0);
 in96 : in unsigned(7 downto 0);
 in97 : in unsigned(7 downto 0);
 in98 : in unsigned(7 downto 0);
 in99 : in unsigned(7 downto 0);
 in100 : in unsigned(7 downto 0);
 in101 : in unsigned(7 downto 0);
 in102 : in unsigned(7 downto 0);
 in103 : in unsigned(7 downto 0);
 in104 : in unsigned(7 downto 0);
 in105 : in unsigned(7 downto 0);
 in106 : in unsigned(7 downto 0);
 in107 : in unsigned(7 downto 0);
 in108 : in unsigned(7 downto 0);
 in109 : in unsigned(7 downto 0);
 in110 : in unsigned(7 downto 0);
 in111 : in unsigned(7 downto 0);
 in112 : in unsigned(7 downto 0);
 in113 : in unsigned(7 downto 0);
 in114 : in unsigned(7 downto 0);
 in115 : in unsigned(7 downto 0);
 in116 : in unsigned(7 downto 0);
 in117 : in unsigned(7 downto 0);
 in118 : in unsigned(7 downto 0);
 in119 : in unsigned(7 downto 0);
 in120 : in unsigned(7 downto 0);
 in121 : in unsigned(7 downto 0);
 in122 : in unsigned(7 downto 0);
 in123 : in unsigned(7 downto 0);
 in124 : in unsigned(7 downto 0);
 in125 : in unsigned(7 downto 0);
 in126 : in unsigned(7 downto 0);
 in127 : in unsigned(7 downto 0);
 return_output : out unsigned(7 downto 0));
end uint8_mux128_0CLK_9347d63d;
architecture arch of uint8_mux128_0CLK_9347d63d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_85c1]
signal layer0_node0_MUX_bit_math_h_l18_c3_85c1_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_85c1_iftrue : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_85c1_iffalse : unsigned(7 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_85c1_return_output : unsigned(7 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_a7d4]
signal layer0_node1_MUX_bit_math_h_l29_c3_a7d4_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iftrue : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iffalse : unsigned(7 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_a7d4_return_output : unsigned(7 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_43b7]
signal layer0_node2_MUX_bit_math_h_l40_c3_43b7_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_43b7_iftrue : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_43b7_iffalse : unsigned(7 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_43b7_return_output : unsigned(7 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_a274]
signal layer0_node3_MUX_bit_math_h_l51_c3_a274_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_a274_iftrue : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_a274_iffalse : unsigned(7 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_a274_return_output : unsigned(7 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_2eec]
signal layer0_node4_MUX_bit_math_h_l62_c3_2eec_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_2eec_iftrue : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_2eec_iffalse : unsigned(7 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_2eec_return_output : unsigned(7 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_5736]
signal layer0_node5_MUX_bit_math_h_l73_c3_5736_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_5736_iftrue : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_5736_iffalse : unsigned(7 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_5736_return_output : unsigned(7 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_62aa]
signal layer0_node6_MUX_bit_math_h_l84_c3_62aa_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_62aa_iftrue : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_62aa_iffalse : unsigned(7 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_62aa_return_output : unsigned(7 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_c2e4]
signal layer0_node7_MUX_bit_math_h_l95_c3_c2e4_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iftrue : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iffalse : unsigned(7 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_c2e4_return_output : unsigned(7 downto 0);

-- layer0_node8_MUX[bit_math_h_l106_c3_22f1]
signal layer0_node8_MUX_bit_math_h_l106_c3_22f1_cond : unsigned(0 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_22f1_iftrue : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_22f1_iffalse : unsigned(7 downto 0);
signal layer0_node8_MUX_bit_math_h_l106_c3_22f1_return_output : unsigned(7 downto 0);

-- layer0_node9_MUX[bit_math_h_l117_c3_391b]
signal layer0_node9_MUX_bit_math_h_l117_c3_391b_cond : unsigned(0 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_391b_iftrue : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_391b_iffalse : unsigned(7 downto 0);
signal layer0_node9_MUX_bit_math_h_l117_c3_391b_return_output : unsigned(7 downto 0);

-- layer0_node10_MUX[bit_math_h_l128_c3_1e58]
signal layer0_node10_MUX_bit_math_h_l128_c3_1e58_cond : unsigned(0 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_1e58_iftrue : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_1e58_iffalse : unsigned(7 downto 0);
signal layer0_node10_MUX_bit_math_h_l128_c3_1e58_return_output : unsigned(7 downto 0);

-- layer0_node11_MUX[bit_math_h_l139_c3_6d2d]
signal layer0_node11_MUX_bit_math_h_l139_c3_6d2d_cond : unsigned(0 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iftrue : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iffalse : unsigned(7 downto 0);
signal layer0_node11_MUX_bit_math_h_l139_c3_6d2d_return_output : unsigned(7 downto 0);

-- layer0_node12_MUX[bit_math_h_l150_c3_40e1]
signal layer0_node12_MUX_bit_math_h_l150_c3_40e1_cond : unsigned(0 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_40e1_iftrue : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_40e1_iffalse : unsigned(7 downto 0);
signal layer0_node12_MUX_bit_math_h_l150_c3_40e1_return_output : unsigned(7 downto 0);

-- layer0_node13_MUX[bit_math_h_l161_c3_28f7]
signal layer0_node13_MUX_bit_math_h_l161_c3_28f7_cond : unsigned(0 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_28f7_iftrue : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_28f7_iffalse : unsigned(7 downto 0);
signal layer0_node13_MUX_bit_math_h_l161_c3_28f7_return_output : unsigned(7 downto 0);

-- layer0_node14_MUX[bit_math_h_l172_c3_e31d]
signal layer0_node14_MUX_bit_math_h_l172_c3_e31d_cond : unsigned(0 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_e31d_iftrue : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_e31d_iffalse : unsigned(7 downto 0);
signal layer0_node14_MUX_bit_math_h_l172_c3_e31d_return_output : unsigned(7 downto 0);

-- layer0_node15_MUX[bit_math_h_l183_c3_313e]
signal layer0_node15_MUX_bit_math_h_l183_c3_313e_cond : unsigned(0 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_313e_iftrue : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_313e_iffalse : unsigned(7 downto 0);
signal layer0_node15_MUX_bit_math_h_l183_c3_313e_return_output : unsigned(7 downto 0);

-- layer0_node16_MUX[bit_math_h_l194_c3_614a]
signal layer0_node16_MUX_bit_math_h_l194_c3_614a_cond : unsigned(0 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_614a_iftrue : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_614a_iffalse : unsigned(7 downto 0);
signal layer0_node16_MUX_bit_math_h_l194_c3_614a_return_output : unsigned(7 downto 0);

-- layer0_node17_MUX[bit_math_h_l205_c3_ec06]
signal layer0_node17_MUX_bit_math_h_l205_c3_ec06_cond : unsigned(0 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_ec06_iftrue : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_ec06_iffalse : unsigned(7 downto 0);
signal layer0_node17_MUX_bit_math_h_l205_c3_ec06_return_output : unsigned(7 downto 0);

-- layer0_node18_MUX[bit_math_h_l216_c3_7962]
signal layer0_node18_MUX_bit_math_h_l216_c3_7962_cond : unsigned(0 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_7962_iftrue : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_7962_iffalse : unsigned(7 downto 0);
signal layer0_node18_MUX_bit_math_h_l216_c3_7962_return_output : unsigned(7 downto 0);

-- layer0_node19_MUX[bit_math_h_l227_c3_0da7]
signal layer0_node19_MUX_bit_math_h_l227_c3_0da7_cond : unsigned(0 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_0da7_iftrue : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_0da7_iffalse : unsigned(7 downto 0);
signal layer0_node19_MUX_bit_math_h_l227_c3_0da7_return_output : unsigned(7 downto 0);

-- layer0_node20_MUX[bit_math_h_l238_c3_a0ec]
signal layer0_node20_MUX_bit_math_h_l238_c3_a0ec_cond : unsigned(0 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iftrue : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iffalse : unsigned(7 downto 0);
signal layer0_node20_MUX_bit_math_h_l238_c3_a0ec_return_output : unsigned(7 downto 0);

-- layer0_node21_MUX[bit_math_h_l249_c3_a3f0]
signal layer0_node21_MUX_bit_math_h_l249_c3_a3f0_cond : unsigned(0 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iftrue : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iffalse : unsigned(7 downto 0);
signal layer0_node21_MUX_bit_math_h_l249_c3_a3f0_return_output : unsigned(7 downto 0);

-- layer0_node22_MUX[bit_math_h_l260_c3_50aa]
signal layer0_node22_MUX_bit_math_h_l260_c3_50aa_cond : unsigned(0 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_50aa_iftrue : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_50aa_iffalse : unsigned(7 downto 0);
signal layer0_node22_MUX_bit_math_h_l260_c3_50aa_return_output : unsigned(7 downto 0);

-- layer0_node23_MUX[bit_math_h_l271_c3_b2cd]
signal layer0_node23_MUX_bit_math_h_l271_c3_b2cd_cond : unsigned(0 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iftrue : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iffalse : unsigned(7 downto 0);
signal layer0_node23_MUX_bit_math_h_l271_c3_b2cd_return_output : unsigned(7 downto 0);

-- layer0_node24_MUX[bit_math_h_l282_c3_0847]
signal layer0_node24_MUX_bit_math_h_l282_c3_0847_cond : unsigned(0 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_0847_iftrue : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_0847_iffalse : unsigned(7 downto 0);
signal layer0_node24_MUX_bit_math_h_l282_c3_0847_return_output : unsigned(7 downto 0);

-- layer0_node25_MUX[bit_math_h_l293_c3_d8bb]
signal layer0_node25_MUX_bit_math_h_l293_c3_d8bb_cond : unsigned(0 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iftrue : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iffalse : unsigned(7 downto 0);
signal layer0_node25_MUX_bit_math_h_l293_c3_d8bb_return_output : unsigned(7 downto 0);

-- layer0_node26_MUX[bit_math_h_l304_c3_809a]
signal layer0_node26_MUX_bit_math_h_l304_c3_809a_cond : unsigned(0 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_809a_iftrue : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_809a_iffalse : unsigned(7 downto 0);
signal layer0_node26_MUX_bit_math_h_l304_c3_809a_return_output : unsigned(7 downto 0);

-- layer0_node27_MUX[bit_math_h_l315_c3_a6a8]
signal layer0_node27_MUX_bit_math_h_l315_c3_a6a8_cond : unsigned(0 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iftrue : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iffalse : unsigned(7 downto 0);
signal layer0_node27_MUX_bit_math_h_l315_c3_a6a8_return_output : unsigned(7 downto 0);

-- layer0_node28_MUX[bit_math_h_l326_c3_b62d]
signal layer0_node28_MUX_bit_math_h_l326_c3_b62d_cond : unsigned(0 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_b62d_iftrue : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_b62d_iffalse : unsigned(7 downto 0);
signal layer0_node28_MUX_bit_math_h_l326_c3_b62d_return_output : unsigned(7 downto 0);

-- layer0_node29_MUX[bit_math_h_l337_c3_1d84]
signal layer0_node29_MUX_bit_math_h_l337_c3_1d84_cond : unsigned(0 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_1d84_iftrue : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_1d84_iffalse : unsigned(7 downto 0);
signal layer0_node29_MUX_bit_math_h_l337_c3_1d84_return_output : unsigned(7 downto 0);

-- layer0_node30_MUX[bit_math_h_l348_c3_27f8]
signal layer0_node30_MUX_bit_math_h_l348_c3_27f8_cond : unsigned(0 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_27f8_iftrue : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_27f8_iffalse : unsigned(7 downto 0);
signal layer0_node30_MUX_bit_math_h_l348_c3_27f8_return_output : unsigned(7 downto 0);

-- layer0_node31_MUX[bit_math_h_l359_c3_e962]
signal layer0_node31_MUX_bit_math_h_l359_c3_e962_cond : unsigned(0 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_e962_iftrue : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_e962_iffalse : unsigned(7 downto 0);
signal layer0_node31_MUX_bit_math_h_l359_c3_e962_return_output : unsigned(7 downto 0);

-- layer0_node32_MUX[bit_math_h_l370_c3_45be]
signal layer0_node32_MUX_bit_math_h_l370_c3_45be_cond : unsigned(0 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_45be_iftrue : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_45be_iffalse : unsigned(7 downto 0);
signal layer0_node32_MUX_bit_math_h_l370_c3_45be_return_output : unsigned(7 downto 0);

-- layer0_node33_MUX[bit_math_h_l381_c3_2a50]
signal layer0_node33_MUX_bit_math_h_l381_c3_2a50_cond : unsigned(0 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_2a50_iftrue : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_2a50_iffalse : unsigned(7 downto 0);
signal layer0_node33_MUX_bit_math_h_l381_c3_2a50_return_output : unsigned(7 downto 0);

-- layer0_node34_MUX[bit_math_h_l392_c3_7b48]
signal layer0_node34_MUX_bit_math_h_l392_c3_7b48_cond : unsigned(0 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_7b48_iftrue : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_7b48_iffalse : unsigned(7 downto 0);
signal layer0_node34_MUX_bit_math_h_l392_c3_7b48_return_output : unsigned(7 downto 0);

-- layer0_node35_MUX[bit_math_h_l403_c3_37e5]
signal layer0_node35_MUX_bit_math_h_l403_c3_37e5_cond : unsigned(0 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_37e5_iftrue : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_37e5_iffalse : unsigned(7 downto 0);
signal layer0_node35_MUX_bit_math_h_l403_c3_37e5_return_output : unsigned(7 downto 0);

-- layer0_node36_MUX[bit_math_h_l414_c3_fd1a]
signal layer0_node36_MUX_bit_math_h_l414_c3_fd1a_cond : unsigned(0 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iftrue : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iffalse : unsigned(7 downto 0);
signal layer0_node36_MUX_bit_math_h_l414_c3_fd1a_return_output : unsigned(7 downto 0);

-- layer0_node37_MUX[bit_math_h_l425_c3_8edb]
signal layer0_node37_MUX_bit_math_h_l425_c3_8edb_cond : unsigned(0 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_8edb_iftrue : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_8edb_iffalse : unsigned(7 downto 0);
signal layer0_node37_MUX_bit_math_h_l425_c3_8edb_return_output : unsigned(7 downto 0);

-- layer0_node38_MUX[bit_math_h_l436_c3_b87e]
signal layer0_node38_MUX_bit_math_h_l436_c3_b87e_cond : unsigned(0 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_b87e_iftrue : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_b87e_iffalse : unsigned(7 downto 0);
signal layer0_node38_MUX_bit_math_h_l436_c3_b87e_return_output : unsigned(7 downto 0);

-- layer0_node39_MUX[bit_math_h_l447_c3_8780]
signal layer0_node39_MUX_bit_math_h_l447_c3_8780_cond : unsigned(0 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_8780_iftrue : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_8780_iffalse : unsigned(7 downto 0);
signal layer0_node39_MUX_bit_math_h_l447_c3_8780_return_output : unsigned(7 downto 0);

-- layer0_node40_MUX[bit_math_h_l458_c3_a82d]
signal layer0_node40_MUX_bit_math_h_l458_c3_a82d_cond : unsigned(0 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_a82d_iftrue : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_a82d_iffalse : unsigned(7 downto 0);
signal layer0_node40_MUX_bit_math_h_l458_c3_a82d_return_output : unsigned(7 downto 0);

-- layer0_node41_MUX[bit_math_h_l469_c3_f332]
signal layer0_node41_MUX_bit_math_h_l469_c3_f332_cond : unsigned(0 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_f332_iftrue : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_f332_iffalse : unsigned(7 downto 0);
signal layer0_node41_MUX_bit_math_h_l469_c3_f332_return_output : unsigned(7 downto 0);

-- layer0_node42_MUX[bit_math_h_l480_c3_8296]
signal layer0_node42_MUX_bit_math_h_l480_c3_8296_cond : unsigned(0 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_8296_iftrue : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_8296_iffalse : unsigned(7 downto 0);
signal layer0_node42_MUX_bit_math_h_l480_c3_8296_return_output : unsigned(7 downto 0);

-- layer0_node43_MUX[bit_math_h_l491_c3_a5e9]
signal layer0_node43_MUX_bit_math_h_l491_c3_a5e9_cond : unsigned(0 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iftrue : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iffalse : unsigned(7 downto 0);
signal layer0_node43_MUX_bit_math_h_l491_c3_a5e9_return_output : unsigned(7 downto 0);

-- layer0_node44_MUX[bit_math_h_l502_c3_7ff6]
signal layer0_node44_MUX_bit_math_h_l502_c3_7ff6_cond : unsigned(0 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iftrue : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iffalse : unsigned(7 downto 0);
signal layer0_node44_MUX_bit_math_h_l502_c3_7ff6_return_output : unsigned(7 downto 0);

-- layer0_node45_MUX[bit_math_h_l513_c3_1806]
signal layer0_node45_MUX_bit_math_h_l513_c3_1806_cond : unsigned(0 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_1806_iftrue : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_1806_iffalse : unsigned(7 downto 0);
signal layer0_node45_MUX_bit_math_h_l513_c3_1806_return_output : unsigned(7 downto 0);

-- layer0_node46_MUX[bit_math_h_l524_c3_c07c]
signal layer0_node46_MUX_bit_math_h_l524_c3_c07c_cond : unsigned(0 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_c07c_iftrue : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_c07c_iffalse : unsigned(7 downto 0);
signal layer0_node46_MUX_bit_math_h_l524_c3_c07c_return_output : unsigned(7 downto 0);

-- layer0_node47_MUX[bit_math_h_l535_c3_a2fb]
signal layer0_node47_MUX_bit_math_h_l535_c3_a2fb_cond : unsigned(0 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iftrue : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iffalse : unsigned(7 downto 0);
signal layer0_node47_MUX_bit_math_h_l535_c3_a2fb_return_output : unsigned(7 downto 0);

-- layer0_node48_MUX[bit_math_h_l546_c3_a700]
signal layer0_node48_MUX_bit_math_h_l546_c3_a700_cond : unsigned(0 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_a700_iftrue : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_a700_iffalse : unsigned(7 downto 0);
signal layer0_node48_MUX_bit_math_h_l546_c3_a700_return_output : unsigned(7 downto 0);

-- layer0_node49_MUX[bit_math_h_l557_c3_5e53]
signal layer0_node49_MUX_bit_math_h_l557_c3_5e53_cond : unsigned(0 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_5e53_iftrue : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_5e53_iffalse : unsigned(7 downto 0);
signal layer0_node49_MUX_bit_math_h_l557_c3_5e53_return_output : unsigned(7 downto 0);

-- layer0_node50_MUX[bit_math_h_l568_c3_ac6c]
signal layer0_node50_MUX_bit_math_h_l568_c3_ac6c_cond : unsigned(0 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iftrue : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iffalse : unsigned(7 downto 0);
signal layer0_node50_MUX_bit_math_h_l568_c3_ac6c_return_output : unsigned(7 downto 0);

-- layer0_node51_MUX[bit_math_h_l579_c3_c608]
signal layer0_node51_MUX_bit_math_h_l579_c3_c608_cond : unsigned(0 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_c608_iftrue : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_c608_iffalse : unsigned(7 downto 0);
signal layer0_node51_MUX_bit_math_h_l579_c3_c608_return_output : unsigned(7 downto 0);

-- layer0_node52_MUX[bit_math_h_l590_c3_f975]
signal layer0_node52_MUX_bit_math_h_l590_c3_f975_cond : unsigned(0 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_f975_iftrue : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_f975_iffalse : unsigned(7 downto 0);
signal layer0_node52_MUX_bit_math_h_l590_c3_f975_return_output : unsigned(7 downto 0);

-- layer0_node53_MUX[bit_math_h_l601_c3_86a8]
signal layer0_node53_MUX_bit_math_h_l601_c3_86a8_cond : unsigned(0 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_86a8_iftrue : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_86a8_iffalse : unsigned(7 downto 0);
signal layer0_node53_MUX_bit_math_h_l601_c3_86a8_return_output : unsigned(7 downto 0);

-- layer0_node54_MUX[bit_math_h_l612_c3_21f7]
signal layer0_node54_MUX_bit_math_h_l612_c3_21f7_cond : unsigned(0 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_21f7_iftrue : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_21f7_iffalse : unsigned(7 downto 0);
signal layer0_node54_MUX_bit_math_h_l612_c3_21f7_return_output : unsigned(7 downto 0);

-- layer0_node55_MUX[bit_math_h_l623_c3_a654]
signal layer0_node55_MUX_bit_math_h_l623_c3_a654_cond : unsigned(0 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_a654_iftrue : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_a654_iffalse : unsigned(7 downto 0);
signal layer0_node55_MUX_bit_math_h_l623_c3_a654_return_output : unsigned(7 downto 0);

-- layer0_node56_MUX[bit_math_h_l634_c3_259e]
signal layer0_node56_MUX_bit_math_h_l634_c3_259e_cond : unsigned(0 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_259e_iftrue : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_259e_iffalse : unsigned(7 downto 0);
signal layer0_node56_MUX_bit_math_h_l634_c3_259e_return_output : unsigned(7 downto 0);

-- layer0_node57_MUX[bit_math_h_l645_c3_3acf]
signal layer0_node57_MUX_bit_math_h_l645_c3_3acf_cond : unsigned(0 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_3acf_iftrue : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_3acf_iffalse : unsigned(7 downto 0);
signal layer0_node57_MUX_bit_math_h_l645_c3_3acf_return_output : unsigned(7 downto 0);

-- layer0_node58_MUX[bit_math_h_l656_c3_6a0d]
signal layer0_node58_MUX_bit_math_h_l656_c3_6a0d_cond : unsigned(0 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iftrue : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iffalse : unsigned(7 downto 0);
signal layer0_node58_MUX_bit_math_h_l656_c3_6a0d_return_output : unsigned(7 downto 0);

-- layer0_node59_MUX[bit_math_h_l667_c3_060a]
signal layer0_node59_MUX_bit_math_h_l667_c3_060a_cond : unsigned(0 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_060a_iftrue : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_060a_iffalse : unsigned(7 downto 0);
signal layer0_node59_MUX_bit_math_h_l667_c3_060a_return_output : unsigned(7 downto 0);

-- layer0_node60_MUX[bit_math_h_l678_c3_dedf]
signal layer0_node60_MUX_bit_math_h_l678_c3_dedf_cond : unsigned(0 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_dedf_iftrue : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_dedf_iffalse : unsigned(7 downto 0);
signal layer0_node60_MUX_bit_math_h_l678_c3_dedf_return_output : unsigned(7 downto 0);

-- layer0_node61_MUX[bit_math_h_l689_c3_26a3]
signal layer0_node61_MUX_bit_math_h_l689_c3_26a3_cond : unsigned(0 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_26a3_iftrue : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_26a3_iffalse : unsigned(7 downto 0);
signal layer0_node61_MUX_bit_math_h_l689_c3_26a3_return_output : unsigned(7 downto 0);

-- layer0_node62_MUX[bit_math_h_l700_c3_7046]
signal layer0_node62_MUX_bit_math_h_l700_c3_7046_cond : unsigned(0 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_7046_iftrue : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_7046_iffalse : unsigned(7 downto 0);
signal layer0_node62_MUX_bit_math_h_l700_c3_7046_return_output : unsigned(7 downto 0);

-- layer0_node63_MUX[bit_math_h_l711_c3_0125]
signal layer0_node63_MUX_bit_math_h_l711_c3_0125_cond : unsigned(0 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_0125_iftrue : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_0125_iffalse : unsigned(7 downto 0);
signal layer0_node63_MUX_bit_math_h_l711_c3_0125_return_output : unsigned(7 downto 0);

-- layer1_node0_MUX[bit_math_h_l728_c3_287e]
signal layer1_node0_MUX_bit_math_h_l728_c3_287e_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_287e_iftrue : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_287e_iffalse : unsigned(7 downto 0);
signal layer1_node0_MUX_bit_math_h_l728_c3_287e_return_output : unsigned(7 downto 0);

-- layer1_node1_MUX[bit_math_h_l739_c3_3eb3]
signal layer1_node1_MUX_bit_math_h_l739_c3_3eb3_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iftrue : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iffalse : unsigned(7 downto 0);
signal layer1_node1_MUX_bit_math_h_l739_c3_3eb3_return_output : unsigned(7 downto 0);

-- layer1_node2_MUX[bit_math_h_l750_c3_e4a0]
signal layer1_node2_MUX_bit_math_h_l750_c3_e4a0_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iftrue : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iffalse : unsigned(7 downto 0);
signal layer1_node2_MUX_bit_math_h_l750_c3_e4a0_return_output : unsigned(7 downto 0);

-- layer1_node3_MUX[bit_math_h_l761_c3_123f]
signal layer1_node3_MUX_bit_math_h_l761_c3_123f_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_123f_iftrue : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_123f_iffalse : unsigned(7 downto 0);
signal layer1_node3_MUX_bit_math_h_l761_c3_123f_return_output : unsigned(7 downto 0);

-- layer1_node4_MUX[bit_math_h_l772_c3_0289]
signal layer1_node4_MUX_bit_math_h_l772_c3_0289_cond : unsigned(0 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_0289_iftrue : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_0289_iffalse : unsigned(7 downto 0);
signal layer1_node4_MUX_bit_math_h_l772_c3_0289_return_output : unsigned(7 downto 0);

-- layer1_node5_MUX[bit_math_h_l783_c3_58a8]
signal layer1_node5_MUX_bit_math_h_l783_c3_58a8_cond : unsigned(0 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_58a8_iftrue : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_58a8_iffalse : unsigned(7 downto 0);
signal layer1_node5_MUX_bit_math_h_l783_c3_58a8_return_output : unsigned(7 downto 0);

-- layer1_node6_MUX[bit_math_h_l794_c3_ebf4]
signal layer1_node6_MUX_bit_math_h_l794_c3_ebf4_cond : unsigned(0 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iftrue : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iffalse : unsigned(7 downto 0);
signal layer1_node6_MUX_bit_math_h_l794_c3_ebf4_return_output : unsigned(7 downto 0);

-- layer1_node7_MUX[bit_math_h_l805_c3_1224]
signal layer1_node7_MUX_bit_math_h_l805_c3_1224_cond : unsigned(0 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_1224_iftrue : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_1224_iffalse : unsigned(7 downto 0);
signal layer1_node7_MUX_bit_math_h_l805_c3_1224_return_output : unsigned(7 downto 0);

-- layer1_node8_MUX[bit_math_h_l816_c3_db42]
signal layer1_node8_MUX_bit_math_h_l816_c3_db42_cond : unsigned(0 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_db42_iftrue : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_db42_iffalse : unsigned(7 downto 0);
signal layer1_node8_MUX_bit_math_h_l816_c3_db42_return_output : unsigned(7 downto 0);

-- layer1_node9_MUX[bit_math_h_l827_c3_8290]
signal layer1_node9_MUX_bit_math_h_l827_c3_8290_cond : unsigned(0 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_8290_iftrue : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_8290_iffalse : unsigned(7 downto 0);
signal layer1_node9_MUX_bit_math_h_l827_c3_8290_return_output : unsigned(7 downto 0);

-- layer1_node10_MUX[bit_math_h_l838_c3_a2e2]
signal layer1_node10_MUX_bit_math_h_l838_c3_a2e2_cond : unsigned(0 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iftrue : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iffalse : unsigned(7 downto 0);
signal layer1_node10_MUX_bit_math_h_l838_c3_a2e2_return_output : unsigned(7 downto 0);

-- layer1_node11_MUX[bit_math_h_l849_c3_dc54]
signal layer1_node11_MUX_bit_math_h_l849_c3_dc54_cond : unsigned(0 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_dc54_iftrue : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_dc54_iffalse : unsigned(7 downto 0);
signal layer1_node11_MUX_bit_math_h_l849_c3_dc54_return_output : unsigned(7 downto 0);

-- layer1_node12_MUX[bit_math_h_l860_c3_7af8]
signal layer1_node12_MUX_bit_math_h_l860_c3_7af8_cond : unsigned(0 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_7af8_iftrue : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_7af8_iffalse : unsigned(7 downto 0);
signal layer1_node12_MUX_bit_math_h_l860_c3_7af8_return_output : unsigned(7 downto 0);

-- layer1_node13_MUX[bit_math_h_l871_c3_d1fd]
signal layer1_node13_MUX_bit_math_h_l871_c3_d1fd_cond : unsigned(0 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iftrue : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iffalse : unsigned(7 downto 0);
signal layer1_node13_MUX_bit_math_h_l871_c3_d1fd_return_output : unsigned(7 downto 0);

-- layer1_node14_MUX[bit_math_h_l882_c3_10cf]
signal layer1_node14_MUX_bit_math_h_l882_c3_10cf_cond : unsigned(0 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_10cf_iftrue : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_10cf_iffalse : unsigned(7 downto 0);
signal layer1_node14_MUX_bit_math_h_l882_c3_10cf_return_output : unsigned(7 downto 0);

-- layer1_node15_MUX[bit_math_h_l893_c3_3f51]
signal layer1_node15_MUX_bit_math_h_l893_c3_3f51_cond : unsigned(0 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_3f51_iftrue : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_3f51_iffalse : unsigned(7 downto 0);
signal layer1_node15_MUX_bit_math_h_l893_c3_3f51_return_output : unsigned(7 downto 0);

-- layer1_node16_MUX[bit_math_h_l904_c3_e9a5]
signal layer1_node16_MUX_bit_math_h_l904_c3_e9a5_cond : unsigned(0 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iftrue : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iffalse : unsigned(7 downto 0);
signal layer1_node16_MUX_bit_math_h_l904_c3_e9a5_return_output : unsigned(7 downto 0);

-- layer1_node17_MUX[bit_math_h_l915_c3_4b4e]
signal layer1_node17_MUX_bit_math_h_l915_c3_4b4e_cond : unsigned(0 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iftrue : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iffalse : unsigned(7 downto 0);
signal layer1_node17_MUX_bit_math_h_l915_c3_4b4e_return_output : unsigned(7 downto 0);

-- layer1_node18_MUX[bit_math_h_l926_c3_5844]
signal layer1_node18_MUX_bit_math_h_l926_c3_5844_cond : unsigned(0 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_5844_iftrue : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_5844_iffalse : unsigned(7 downto 0);
signal layer1_node18_MUX_bit_math_h_l926_c3_5844_return_output : unsigned(7 downto 0);

-- layer1_node19_MUX[bit_math_h_l937_c3_7dba]
signal layer1_node19_MUX_bit_math_h_l937_c3_7dba_cond : unsigned(0 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_7dba_iftrue : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_7dba_iffalse : unsigned(7 downto 0);
signal layer1_node19_MUX_bit_math_h_l937_c3_7dba_return_output : unsigned(7 downto 0);

-- layer1_node20_MUX[bit_math_h_l948_c3_2725]
signal layer1_node20_MUX_bit_math_h_l948_c3_2725_cond : unsigned(0 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2725_iftrue : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2725_iffalse : unsigned(7 downto 0);
signal layer1_node20_MUX_bit_math_h_l948_c3_2725_return_output : unsigned(7 downto 0);

-- layer1_node21_MUX[bit_math_h_l959_c3_8499]
signal layer1_node21_MUX_bit_math_h_l959_c3_8499_cond : unsigned(0 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_8499_iftrue : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_8499_iffalse : unsigned(7 downto 0);
signal layer1_node21_MUX_bit_math_h_l959_c3_8499_return_output : unsigned(7 downto 0);

-- layer1_node22_MUX[bit_math_h_l970_c3_65bd]
signal layer1_node22_MUX_bit_math_h_l970_c3_65bd_cond : unsigned(0 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_65bd_iftrue : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_65bd_iffalse : unsigned(7 downto 0);
signal layer1_node22_MUX_bit_math_h_l970_c3_65bd_return_output : unsigned(7 downto 0);

-- layer1_node23_MUX[bit_math_h_l981_c3_3335]
signal layer1_node23_MUX_bit_math_h_l981_c3_3335_cond : unsigned(0 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_3335_iftrue : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_3335_iffalse : unsigned(7 downto 0);
signal layer1_node23_MUX_bit_math_h_l981_c3_3335_return_output : unsigned(7 downto 0);

-- layer1_node24_MUX[bit_math_h_l992_c3_8ee7]
signal layer1_node24_MUX_bit_math_h_l992_c3_8ee7_cond : unsigned(0 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iftrue : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iffalse : unsigned(7 downto 0);
signal layer1_node24_MUX_bit_math_h_l992_c3_8ee7_return_output : unsigned(7 downto 0);

-- layer1_node25_MUX[bit_math_h_l1003_c3_8e94]
signal layer1_node25_MUX_bit_math_h_l1003_c3_8e94_cond : unsigned(0 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iftrue : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iffalse : unsigned(7 downto 0);
signal layer1_node25_MUX_bit_math_h_l1003_c3_8e94_return_output : unsigned(7 downto 0);

-- layer1_node26_MUX[bit_math_h_l1014_c3_d8aa]
signal layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_cond : unsigned(0 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iftrue : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iffalse : unsigned(7 downto 0);
signal layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_return_output : unsigned(7 downto 0);

-- layer1_node27_MUX[bit_math_h_l1025_c3_465f]
signal layer1_node27_MUX_bit_math_h_l1025_c3_465f_cond : unsigned(0 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_465f_iftrue : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_465f_iffalse : unsigned(7 downto 0);
signal layer1_node27_MUX_bit_math_h_l1025_c3_465f_return_output : unsigned(7 downto 0);

-- layer1_node28_MUX[bit_math_h_l1036_c3_f568]
signal layer1_node28_MUX_bit_math_h_l1036_c3_f568_cond : unsigned(0 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_f568_iftrue : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_f568_iffalse : unsigned(7 downto 0);
signal layer1_node28_MUX_bit_math_h_l1036_c3_f568_return_output : unsigned(7 downto 0);

-- layer1_node29_MUX[bit_math_h_l1047_c3_8f77]
signal layer1_node29_MUX_bit_math_h_l1047_c3_8f77_cond : unsigned(0 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iftrue : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iffalse : unsigned(7 downto 0);
signal layer1_node29_MUX_bit_math_h_l1047_c3_8f77_return_output : unsigned(7 downto 0);

-- layer1_node30_MUX[bit_math_h_l1058_c3_d4dc]
signal layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_cond : unsigned(0 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iftrue : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iffalse : unsigned(7 downto 0);
signal layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_return_output : unsigned(7 downto 0);

-- layer1_node31_MUX[bit_math_h_l1069_c3_6881]
signal layer1_node31_MUX_bit_math_h_l1069_c3_6881_cond : unsigned(0 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_6881_iftrue : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_6881_iffalse : unsigned(7 downto 0);
signal layer1_node31_MUX_bit_math_h_l1069_c3_6881_return_output : unsigned(7 downto 0);

-- layer2_node0_MUX[bit_math_h_l1086_c3_f1d8]
signal layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iftrue : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iffalse : unsigned(7 downto 0);
signal layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_return_output : unsigned(7 downto 0);

-- layer2_node1_MUX[bit_math_h_l1097_c3_1a30]
signal layer2_node1_MUX_bit_math_h_l1097_c3_1a30_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iftrue : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iffalse : unsigned(7 downto 0);
signal layer2_node1_MUX_bit_math_h_l1097_c3_1a30_return_output : unsigned(7 downto 0);

-- layer2_node2_MUX[bit_math_h_l1108_c3_0b56]
signal layer2_node2_MUX_bit_math_h_l1108_c3_0b56_cond : unsigned(0 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iftrue : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iffalse : unsigned(7 downto 0);
signal layer2_node2_MUX_bit_math_h_l1108_c3_0b56_return_output : unsigned(7 downto 0);

-- layer2_node3_MUX[bit_math_h_l1119_c3_7df6]
signal layer2_node3_MUX_bit_math_h_l1119_c3_7df6_cond : unsigned(0 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iftrue : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iffalse : unsigned(7 downto 0);
signal layer2_node3_MUX_bit_math_h_l1119_c3_7df6_return_output : unsigned(7 downto 0);

-- layer2_node4_MUX[bit_math_h_l1130_c3_7e5b]
signal layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_cond : unsigned(0 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iftrue : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iffalse : unsigned(7 downto 0);
signal layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_return_output : unsigned(7 downto 0);

-- layer2_node5_MUX[bit_math_h_l1141_c3_25de]
signal layer2_node5_MUX_bit_math_h_l1141_c3_25de_cond : unsigned(0 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_25de_iftrue : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_25de_iffalse : unsigned(7 downto 0);
signal layer2_node5_MUX_bit_math_h_l1141_c3_25de_return_output : unsigned(7 downto 0);

-- layer2_node6_MUX[bit_math_h_l1152_c3_be62]
signal layer2_node6_MUX_bit_math_h_l1152_c3_be62_cond : unsigned(0 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_be62_iftrue : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_be62_iffalse : unsigned(7 downto 0);
signal layer2_node6_MUX_bit_math_h_l1152_c3_be62_return_output : unsigned(7 downto 0);

-- layer2_node7_MUX[bit_math_h_l1163_c3_9403]
signal layer2_node7_MUX_bit_math_h_l1163_c3_9403_cond : unsigned(0 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_9403_iftrue : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_9403_iffalse : unsigned(7 downto 0);
signal layer2_node7_MUX_bit_math_h_l1163_c3_9403_return_output : unsigned(7 downto 0);

-- layer2_node8_MUX[bit_math_h_l1174_c3_918c]
signal layer2_node8_MUX_bit_math_h_l1174_c3_918c_cond : unsigned(0 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_918c_iftrue : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_918c_iffalse : unsigned(7 downto 0);
signal layer2_node8_MUX_bit_math_h_l1174_c3_918c_return_output : unsigned(7 downto 0);

-- layer2_node9_MUX[bit_math_h_l1185_c3_9e4b]
signal layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_cond : unsigned(0 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iftrue : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iffalse : unsigned(7 downto 0);
signal layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_return_output : unsigned(7 downto 0);

-- layer2_node10_MUX[bit_math_h_l1196_c3_3974]
signal layer2_node10_MUX_bit_math_h_l1196_c3_3974_cond : unsigned(0 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_3974_iftrue : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_3974_iffalse : unsigned(7 downto 0);
signal layer2_node10_MUX_bit_math_h_l1196_c3_3974_return_output : unsigned(7 downto 0);

-- layer2_node11_MUX[bit_math_h_l1207_c3_80d7]
signal layer2_node11_MUX_bit_math_h_l1207_c3_80d7_cond : unsigned(0 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iftrue : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iffalse : unsigned(7 downto 0);
signal layer2_node11_MUX_bit_math_h_l1207_c3_80d7_return_output : unsigned(7 downto 0);

-- layer2_node12_MUX[bit_math_h_l1218_c3_fc60]
signal layer2_node12_MUX_bit_math_h_l1218_c3_fc60_cond : unsigned(0 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iftrue : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iffalse : unsigned(7 downto 0);
signal layer2_node12_MUX_bit_math_h_l1218_c3_fc60_return_output : unsigned(7 downto 0);

-- layer2_node13_MUX[bit_math_h_l1229_c3_6c25]
signal layer2_node13_MUX_bit_math_h_l1229_c3_6c25_cond : unsigned(0 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iftrue : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iffalse : unsigned(7 downto 0);
signal layer2_node13_MUX_bit_math_h_l1229_c3_6c25_return_output : unsigned(7 downto 0);

-- layer2_node14_MUX[bit_math_h_l1240_c3_75b9]
signal layer2_node14_MUX_bit_math_h_l1240_c3_75b9_cond : unsigned(0 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iftrue : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iffalse : unsigned(7 downto 0);
signal layer2_node14_MUX_bit_math_h_l1240_c3_75b9_return_output : unsigned(7 downto 0);

-- layer2_node15_MUX[bit_math_h_l1251_c3_ecd2]
signal layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_cond : unsigned(0 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iftrue : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iffalse : unsigned(7 downto 0);
signal layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_return_output : unsigned(7 downto 0);

-- layer3_node0_MUX[bit_math_h_l1268_c3_324b]
signal layer3_node0_MUX_bit_math_h_l1268_c3_324b_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_324b_iftrue : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_324b_iffalse : unsigned(7 downto 0);
signal layer3_node0_MUX_bit_math_h_l1268_c3_324b_return_output : unsigned(7 downto 0);

-- layer3_node1_MUX[bit_math_h_l1279_c3_eea1]
signal layer3_node1_MUX_bit_math_h_l1279_c3_eea1_cond : unsigned(0 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iftrue : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iffalse : unsigned(7 downto 0);
signal layer3_node1_MUX_bit_math_h_l1279_c3_eea1_return_output : unsigned(7 downto 0);

-- layer3_node2_MUX[bit_math_h_l1290_c3_c56d]
signal layer3_node2_MUX_bit_math_h_l1290_c3_c56d_cond : unsigned(0 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iftrue : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iffalse : unsigned(7 downto 0);
signal layer3_node2_MUX_bit_math_h_l1290_c3_c56d_return_output : unsigned(7 downto 0);

-- layer3_node3_MUX[bit_math_h_l1301_c3_98b1]
signal layer3_node3_MUX_bit_math_h_l1301_c3_98b1_cond : unsigned(0 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iftrue : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iffalse : unsigned(7 downto 0);
signal layer3_node3_MUX_bit_math_h_l1301_c3_98b1_return_output : unsigned(7 downto 0);

-- layer3_node4_MUX[bit_math_h_l1312_c3_4b99]
signal layer3_node4_MUX_bit_math_h_l1312_c3_4b99_cond : unsigned(0 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iftrue : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iffalse : unsigned(7 downto 0);
signal layer3_node4_MUX_bit_math_h_l1312_c3_4b99_return_output : unsigned(7 downto 0);

-- layer3_node5_MUX[bit_math_h_l1323_c3_75a2]
signal layer3_node5_MUX_bit_math_h_l1323_c3_75a2_cond : unsigned(0 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iftrue : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iffalse : unsigned(7 downto 0);
signal layer3_node5_MUX_bit_math_h_l1323_c3_75a2_return_output : unsigned(7 downto 0);

-- layer3_node6_MUX[bit_math_h_l1334_c3_483e]
signal layer3_node6_MUX_bit_math_h_l1334_c3_483e_cond : unsigned(0 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_483e_iftrue : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_483e_iffalse : unsigned(7 downto 0);
signal layer3_node6_MUX_bit_math_h_l1334_c3_483e_return_output : unsigned(7 downto 0);

-- layer3_node7_MUX[bit_math_h_l1345_c3_7c85]
signal layer3_node7_MUX_bit_math_h_l1345_c3_7c85_cond : unsigned(0 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iftrue : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iffalse : unsigned(7 downto 0);
signal layer3_node7_MUX_bit_math_h_l1345_c3_7c85_return_output : unsigned(7 downto 0);

-- layer4_node0_MUX[bit_math_h_l1362_c3_bbba]
signal layer4_node0_MUX_bit_math_h_l1362_c3_bbba_cond : unsigned(0 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iftrue : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iffalse : unsigned(7 downto 0);
signal layer4_node0_MUX_bit_math_h_l1362_c3_bbba_return_output : unsigned(7 downto 0);

-- layer4_node1_MUX[bit_math_h_l1373_c3_31df]
signal layer4_node1_MUX_bit_math_h_l1373_c3_31df_cond : unsigned(0 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_31df_iftrue : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_31df_iffalse : unsigned(7 downto 0);
signal layer4_node1_MUX_bit_math_h_l1373_c3_31df_return_output : unsigned(7 downto 0);

-- layer4_node2_MUX[bit_math_h_l1384_c3_d801]
signal layer4_node2_MUX_bit_math_h_l1384_c3_d801_cond : unsigned(0 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_d801_iftrue : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_d801_iffalse : unsigned(7 downto 0);
signal layer4_node2_MUX_bit_math_h_l1384_c3_d801_return_output : unsigned(7 downto 0);

-- layer4_node3_MUX[bit_math_h_l1395_c3_fa88]
signal layer4_node3_MUX_bit_math_h_l1395_c3_fa88_cond : unsigned(0 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iftrue : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iffalse : unsigned(7 downto 0);
signal layer4_node3_MUX_bit_math_h_l1395_c3_fa88_return_output : unsigned(7 downto 0);

-- layer5_node0_MUX[bit_math_h_l1412_c3_ee13]
signal layer5_node0_MUX_bit_math_h_l1412_c3_ee13_cond : unsigned(0 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iftrue : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iffalse : unsigned(7 downto 0);
signal layer5_node0_MUX_bit_math_h_l1412_c3_ee13_return_output : unsigned(7 downto 0);

-- layer5_node1_MUX[bit_math_h_l1423_c3_93d3]
signal layer5_node1_MUX_bit_math_h_l1423_c3_93d3_cond : unsigned(0 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iftrue : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iffalse : unsigned(7 downto 0);
signal layer5_node1_MUX_bit_math_h_l1423_c3_93d3_return_output : unsigned(7 downto 0);

-- layer6_node0_MUX[bit_math_h_l1440_c3_08eb]
signal layer6_node0_MUX_bit_math_h_l1440_c3_08eb_cond : unsigned(0 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iftrue : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iffalse : unsigned(7 downto 0);
signal layer6_node0_MUX_bit_math_h_l1440_c3_08eb_return_output : unsigned(7 downto 0);

function uint7_0_0( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint7_1_1( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint7_2_2( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint7_3_3( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;

function uint7_4_4( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(4- i);
      end loop;
return return_output;
end function;

function uint7_5_5( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(5- i);
      end loop;
return return_output;
end function;

function uint7_6_6( x : unsigned) return unsigned is
--variable x : unsigned(6 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(6- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_85c1
layer0_node0_MUX_bit_math_h_l18_c3_85c1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_85c1_cond,
layer0_node0_MUX_bit_math_h_l18_c3_85c1_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_85c1_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_85c1_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_a7d4
layer0_node1_MUX_bit_math_h_l29_c3_a7d4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_a7d4_cond,
layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_a7d4_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_43b7
layer0_node2_MUX_bit_math_h_l40_c3_43b7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_43b7_cond,
layer0_node2_MUX_bit_math_h_l40_c3_43b7_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_43b7_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_43b7_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_a274
layer0_node3_MUX_bit_math_h_l51_c3_a274 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_a274_cond,
layer0_node3_MUX_bit_math_h_l51_c3_a274_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_a274_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_a274_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_2eec
layer0_node4_MUX_bit_math_h_l62_c3_2eec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_2eec_cond,
layer0_node4_MUX_bit_math_h_l62_c3_2eec_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_2eec_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_2eec_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_5736
layer0_node5_MUX_bit_math_h_l73_c3_5736 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_5736_cond,
layer0_node5_MUX_bit_math_h_l73_c3_5736_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_5736_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_5736_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_62aa
layer0_node6_MUX_bit_math_h_l84_c3_62aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_62aa_cond,
layer0_node6_MUX_bit_math_h_l84_c3_62aa_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_62aa_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_62aa_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_c2e4
layer0_node7_MUX_bit_math_h_l95_c3_c2e4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_c2e4_cond,
layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_c2e4_return_output);

-- layer0_node8_MUX_bit_math_h_l106_c3_22f1
layer0_node8_MUX_bit_math_h_l106_c3_22f1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node8_MUX_bit_math_h_l106_c3_22f1_cond,
layer0_node8_MUX_bit_math_h_l106_c3_22f1_iftrue,
layer0_node8_MUX_bit_math_h_l106_c3_22f1_iffalse,
layer0_node8_MUX_bit_math_h_l106_c3_22f1_return_output);

-- layer0_node9_MUX_bit_math_h_l117_c3_391b
layer0_node9_MUX_bit_math_h_l117_c3_391b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node9_MUX_bit_math_h_l117_c3_391b_cond,
layer0_node9_MUX_bit_math_h_l117_c3_391b_iftrue,
layer0_node9_MUX_bit_math_h_l117_c3_391b_iffalse,
layer0_node9_MUX_bit_math_h_l117_c3_391b_return_output);

-- layer0_node10_MUX_bit_math_h_l128_c3_1e58
layer0_node10_MUX_bit_math_h_l128_c3_1e58 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node10_MUX_bit_math_h_l128_c3_1e58_cond,
layer0_node10_MUX_bit_math_h_l128_c3_1e58_iftrue,
layer0_node10_MUX_bit_math_h_l128_c3_1e58_iffalse,
layer0_node10_MUX_bit_math_h_l128_c3_1e58_return_output);

-- layer0_node11_MUX_bit_math_h_l139_c3_6d2d
layer0_node11_MUX_bit_math_h_l139_c3_6d2d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node11_MUX_bit_math_h_l139_c3_6d2d_cond,
layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iftrue,
layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iffalse,
layer0_node11_MUX_bit_math_h_l139_c3_6d2d_return_output);

-- layer0_node12_MUX_bit_math_h_l150_c3_40e1
layer0_node12_MUX_bit_math_h_l150_c3_40e1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node12_MUX_bit_math_h_l150_c3_40e1_cond,
layer0_node12_MUX_bit_math_h_l150_c3_40e1_iftrue,
layer0_node12_MUX_bit_math_h_l150_c3_40e1_iffalse,
layer0_node12_MUX_bit_math_h_l150_c3_40e1_return_output);

-- layer0_node13_MUX_bit_math_h_l161_c3_28f7
layer0_node13_MUX_bit_math_h_l161_c3_28f7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node13_MUX_bit_math_h_l161_c3_28f7_cond,
layer0_node13_MUX_bit_math_h_l161_c3_28f7_iftrue,
layer0_node13_MUX_bit_math_h_l161_c3_28f7_iffalse,
layer0_node13_MUX_bit_math_h_l161_c3_28f7_return_output);

-- layer0_node14_MUX_bit_math_h_l172_c3_e31d
layer0_node14_MUX_bit_math_h_l172_c3_e31d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node14_MUX_bit_math_h_l172_c3_e31d_cond,
layer0_node14_MUX_bit_math_h_l172_c3_e31d_iftrue,
layer0_node14_MUX_bit_math_h_l172_c3_e31d_iffalse,
layer0_node14_MUX_bit_math_h_l172_c3_e31d_return_output);

-- layer0_node15_MUX_bit_math_h_l183_c3_313e
layer0_node15_MUX_bit_math_h_l183_c3_313e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node15_MUX_bit_math_h_l183_c3_313e_cond,
layer0_node15_MUX_bit_math_h_l183_c3_313e_iftrue,
layer0_node15_MUX_bit_math_h_l183_c3_313e_iffalse,
layer0_node15_MUX_bit_math_h_l183_c3_313e_return_output);

-- layer0_node16_MUX_bit_math_h_l194_c3_614a
layer0_node16_MUX_bit_math_h_l194_c3_614a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node16_MUX_bit_math_h_l194_c3_614a_cond,
layer0_node16_MUX_bit_math_h_l194_c3_614a_iftrue,
layer0_node16_MUX_bit_math_h_l194_c3_614a_iffalse,
layer0_node16_MUX_bit_math_h_l194_c3_614a_return_output);

-- layer0_node17_MUX_bit_math_h_l205_c3_ec06
layer0_node17_MUX_bit_math_h_l205_c3_ec06 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node17_MUX_bit_math_h_l205_c3_ec06_cond,
layer0_node17_MUX_bit_math_h_l205_c3_ec06_iftrue,
layer0_node17_MUX_bit_math_h_l205_c3_ec06_iffalse,
layer0_node17_MUX_bit_math_h_l205_c3_ec06_return_output);

-- layer0_node18_MUX_bit_math_h_l216_c3_7962
layer0_node18_MUX_bit_math_h_l216_c3_7962 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node18_MUX_bit_math_h_l216_c3_7962_cond,
layer0_node18_MUX_bit_math_h_l216_c3_7962_iftrue,
layer0_node18_MUX_bit_math_h_l216_c3_7962_iffalse,
layer0_node18_MUX_bit_math_h_l216_c3_7962_return_output);

-- layer0_node19_MUX_bit_math_h_l227_c3_0da7
layer0_node19_MUX_bit_math_h_l227_c3_0da7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node19_MUX_bit_math_h_l227_c3_0da7_cond,
layer0_node19_MUX_bit_math_h_l227_c3_0da7_iftrue,
layer0_node19_MUX_bit_math_h_l227_c3_0da7_iffalse,
layer0_node19_MUX_bit_math_h_l227_c3_0da7_return_output);

-- layer0_node20_MUX_bit_math_h_l238_c3_a0ec
layer0_node20_MUX_bit_math_h_l238_c3_a0ec : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node20_MUX_bit_math_h_l238_c3_a0ec_cond,
layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iftrue,
layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iffalse,
layer0_node20_MUX_bit_math_h_l238_c3_a0ec_return_output);

-- layer0_node21_MUX_bit_math_h_l249_c3_a3f0
layer0_node21_MUX_bit_math_h_l249_c3_a3f0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node21_MUX_bit_math_h_l249_c3_a3f0_cond,
layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iftrue,
layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iffalse,
layer0_node21_MUX_bit_math_h_l249_c3_a3f0_return_output);

-- layer0_node22_MUX_bit_math_h_l260_c3_50aa
layer0_node22_MUX_bit_math_h_l260_c3_50aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node22_MUX_bit_math_h_l260_c3_50aa_cond,
layer0_node22_MUX_bit_math_h_l260_c3_50aa_iftrue,
layer0_node22_MUX_bit_math_h_l260_c3_50aa_iffalse,
layer0_node22_MUX_bit_math_h_l260_c3_50aa_return_output);

-- layer0_node23_MUX_bit_math_h_l271_c3_b2cd
layer0_node23_MUX_bit_math_h_l271_c3_b2cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node23_MUX_bit_math_h_l271_c3_b2cd_cond,
layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iftrue,
layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iffalse,
layer0_node23_MUX_bit_math_h_l271_c3_b2cd_return_output);

-- layer0_node24_MUX_bit_math_h_l282_c3_0847
layer0_node24_MUX_bit_math_h_l282_c3_0847 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node24_MUX_bit_math_h_l282_c3_0847_cond,
layer0_node24_MUX_bit_math_h_l282_c3_0847_iftrue,
layer0_node24_MUX_bit_math_h_l282_c3_0847_iffalse,
layer0_node24_MUX_bit_math_h_l282_c3_0847_return_output);

-- layer0_node25_MUX_bit_math_h_l293_c3_d8bb
layer0_node25_MUX_bit_math_h_l293_c3_d8bb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node25_MUX_bit_math_h_l293_c3_d8bb_cond,
layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iftrue,
layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iffalse,
layer0_node25_MUX_bit_math_h_l293_c3_d8bb_return_output);

-- layer0_node26_MUX_bit_math_h_l304_c3_809a
layer0_node26_MUX_bit_math_h_l304_c3_809a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node26_MUX_bit_math_h_l304_c3_809a_cond,
layer0_node26_MUX_bit_math_h_l304_c3_809a_iftrue,
layer0_node26_MUX_bit_math_h_l304_c3_809a_iffalse,
layer0_node26_MUX_bit_math_h_l304_c3_809a_return_output);

-- layer0_node27_MUX_bit_math_h_l315_c3_a6a8
layer0_node27_MUX_bit_math_h_l315_c3_a6a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node27_MUX_bit_math_h_l315_c3_a6a8_cond,
layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iftrue,
layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iffalse,
layer0_node27_MUX_bit_math_h_l315_c3_a6a8_return_output);

-- layer0_node28_MUX_bit_math_h_l326_c3_b62d
layer0_node28_MUX_bit_math_h_l326_c3_b62d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node28_MUX_bit_math_h_l326_c3_b62d_cond,
layer0_node28_MUX_bit_math_h_l326_c3_b62d_iftrue,
layer0_node28_MUX_bit_math_h_l326_c3_b62d_iffalse,
layer0_node28_MUX_bit_math_h_l326_c3_b62d_return_output);

-- layer0_node29_MUX_bit_math_h_l337_c3_1d84
layer0_node29_MUX_bit_math_h_l337_c3_1d84 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node29_MUX_bit_math_h_l337_c3_1d84_cond,
layer0_node29_MUX_bit_math_h_l337_c3_1d84_iftrue,
layer0_node29_MUX_bit_math_h_l337_c3_1d84_iffalse,
layer0_node29_MUX_bit_math_h_l337_c3_1d84_return_output);

-- layer0_node30_MUX_bit_math_h_l348_c3_27f8
layer0_node30_MUX_bit_math_h_l348_c3_27f8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node30_MUX_bit_math_h_l348_c3_27f8_cond,
layer0_node30_MUX_bit_math_h_l348_c3_27f8_iftrue,
layer0_node30_MUX_bit_math_h_l348_c3_27f8_iffalse,
layer0_node30_MUX_bit_math_h_l348_c3_27f8_return_output);

-- layer0_node31_MUX_bit_math_h_l359_c3_e962
layer0_node31_MUX_bit_math_h_l359_c3_e962 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node31_MUX_bit_math_h_l359_c3_e962_cond,
layer0_node31_MUX_bit_math_h_l359_c3_e962_iftrue,
layer0_node31_MUX_bit_math_h_l359_c3_e962_iffalse,
layer0_node31_MUX_bit_math_h_l359_c3_e962_return_output);

-- layer0_node32_MUX_bit_math_h_l370_c3_45be
layer0_node32_MUX_bit_math_h_l370_c3_45be : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node32_MUX_bit_math_h_l370_c3_45be_cond,
layer0_node32_MUX_bit_math_h_l370_c3_45be_iftrue,
layer0_node32_MUX_bit_math_h_l370_c3_45be_iffalse,
layer0_node32_MUX_bit_math_h_l370_c3_45be_return_output);

-- layer0_node33_MUX_bit_math_h_l381_c3_2a50
layer0_node33_MUX_bit_math_h_l381_c3_2a50 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node33_MUX_bit_math_h_l381_c3_2a50_cond,
layer0_node33_MUX_bit_math_h_l381_c3_2a50_iftrue,
layer0_node33_MUX_bit_math_h_l381_c3_2a50_iffalse,
layer0_node33_MUX_bit_math_h_l381_c3_2a50_return_output);

-- layer0_node34_MUX_bit_math_h_l392_c3_7b48
layer0_node34_MUX_bit_math_h_l392_c3_7b48 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node34_MUX_bit_math_h_l392_c3_7b48_cond,
layer0_node34_MUX_bit_math_h_l392_c3_7b48_iftrue,
layer0_node34_MUX_bit_math_h_l392_c3_7b48_iffalse,
layer0_node34_MUX_bit_math_h_l392_c3_7b48_return_output);

-- layer0_node35_MUX_bit_math_h_l403_c3_37e5
layer0_node35_MUX_bit_math_h_l403_c3_37e5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node35_MUX_bit_math_h_l403_c3_37e5_cond,
layer0_node35_MUX_bit_math_h_l403_c3_37e5_iftrue,
layer0_node35_MUX_bit_math_h_l403_c3_37e5_iffalse,
layer0_node35_MUX_bit_math_h_l403_c3_37e5_return_output);

-- layer0_node36_MUX_bit_math_h_l414_c3_fd1a
layer0_node36_MUX_bit_math_h_l414_c3_fd1a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node36_MUX_bit_math_h_l414_c3_fd1a_cond,
layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iftrue,
layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iffalse,
layer0_node36_MUX_bit_math_h_l414_c3_fd1a_return_output);

-- layer0_node37_MUX_bit_math_h_l425_c3_8edb
layer0_node37_MUX_bit_math_h_l425_c3_8edb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node37_MUX_bit_math_h_l425_c3_8edb_cond,
layer0_node37_MUX_bit_math_h_l425_c3_8edb_iftrue,
layer0_node37_MUX_bit_math_h_l425_c3_8edb_iffalse,
layer0_node37_MUX_bit_math_h_l425_c3_8edb_return_output);

-- layer0_node38_MUX_bit_math_h_l436_c3_b87e
layer0_node38_MUX_bit_math_h_l436_c3_b87e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node38_MUX_bit_math_h_l436_c3_b87e_cond,
layer0_node38_MUX_bit_math_h_l436_c3_b87e_iftrue,
layer0_node38_MUX_bit_math_h_l436_c3_b87e_iffalse,
layer0_node38_MUX_bit_math_h_l436_c3_b87e_return_output);

-- layer0_node39_MUX_bit_math_h_l447_c3_8780
layer0_node39_MUX_bit_math_h_l447_c3_8780 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node39_MUX_bit_math_h_l447_c3_8780_cond,
layer0_node39_MUX_bit_math_h_l447_c3_8780_iftrue,
layer0_node39_MUX_bit_math_h_l447_c3_8780_iffalse,
layer0_node39_MUX_bit_math_h_l447_c3_8780_return_output);

-- layer0_node40_MUX_bit_math_h_l458_c3_a82d
layer0_node40_MUX_bit_math_h_l458_c3_a82d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node40_MUX_bit_math_h_l458_c3_a82d_cond,
layer0_node40_MUX_bit_math_h_l458_c3_a82d_iftrue,
layer0_node40_MUX_bit_math_h_l458_c3_a82d_iffalse,
layer0_node40_MUX_bit_math_h_l458_c3_a82d_return_output);

-- layer0_node41_MUX_bit_math_h_l469_c3_f332
layer0_node41_MUX_bit_math_h_l469_c3_f332 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node41_MUX_bit_math_h_l469_c3_f332_cond,
layer0_node41_MUX_bit_math_h_l469_c3_f332_iftrue,
layer0_node41_MUX_bit_math_h_l469_c3_f332_iffalse,
layer0_node41_MUX_bit_math_h_l469_c3_f332_return_output);

-- layer0_node42_MUX_bit_math_h_l480_c3_8296
layer0_node42_MUX_bit_math_h_l480_c3_8296 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node42_MUX_bit_math_h_l480_c3_8296_cond,
layer0_node42_MUX_bit_math_h_l480_c3_8296_iftrue,
layer0_node42_MUX_bit_math_h_l480_c3_8296_iffalse,
layer0_node42_MUX_bit_math_h_l480_c3_8296_return_output);

-- layer0_node43_MUX_bit_math_h_l491_c3_a5e9
layer0_node43_MUX_bit_math_h_l491_c3_a5e9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node43_MUX_bit_math_h_l491_c3_a5e9_cond,
layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iftrue,
layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iffalse,
layer0_node43_MUX_bit_math_h_l491_c3_a5e9_return_output);

-- layer0_node44_MUX_bit_math_h_l502_c3_7ff6
layer0_node44_MUX_bit_math_h_l502_c3_7ff6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node44_MUX_bit_math_h_l502_c3_7ff6_cond,
layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iftrue,
layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iffalse,
layer0_node44_MUX_bit_math_h_l502_c3_7ff6_return_output);

-- layer0_node45_MUX_bit_math_h_l513_c3_1806
layer0_node45_MUX_bit_math_h_l513_c3_1806 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node45_MUX_bit_math_h_l513_c3_1806_cond,
layer0_node45_MUX_bit_math_h_l513_c3_1806_iftrue,
layer0_node45_MUX_bit_math_h_l513_c3_1806_iffalse,
layer0_node45_MUX_bit_math_h_l513_c3_1806_return_output);

-- layer0_node46_MUX_bit_math_h_l524_c3_c07c
layer0_node46_MUX_bit_math_h_l524_c3_c07c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node46_MUX_bit_math_h_l524_c3_c07c_cond,
layer0_node46_MUX_bit_math_h_l524_c3_c07c_iftrue,
layer0_node46_MUX_bit_math_h_l524_c3_c07c_iffalse,
layer0_node46_MUX_bit_math_h_l524_c3_c07c_return_output);

-- layer0_node47_MUX_bit_math_h_l535_c3_a2fb
layer0_node47_MUX_bit_math_h_l535_c3_a2fb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node47_MUX_bit_math_h_l535_c3_a2fb_cond,
layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iftrue,
layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iffalse,
layer0_node47_MUX_bit_math_h_l535_c3_a2fb_return_output);

-- layer0_node48_MUX_bit_math_h_l546_c3_a700
layer0_node48_MUX_bit_math_h_l546_c3_a700 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node48_MUX_bit_math_h_l546_c3_a700_cond,
layer0_node48_MUX_bit_math_h_l546_c3_a700_iftrue,
layer0_node48_MUX_bit_math_h_l546_c3_a700_iffalse,
layer0_node48_MUX_bit_math_h_l546_c3_a700_return_output);

-- layer0_node49_MUX_bit_math_h_l557_c3_5e53
layer0_node49_MUX_bit_math_h_l557_c3_5e53 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node49_MUX_bit_math_h_l557_c3_5e53_cond,
layer0_node49_MUX_bit_math_h_l557_c3_5e53_iftrue,
layer0_node49_MUX_bit_math_h_l557_c3_5e53_iffalse,
layer0_node49_MUX_bit_math_h_l557_c3_5e53_return_output);

-- layer0_node50_MUX_bit_math_h_l568_c3_ac6c
layer0_node50_MUX_bit_math_h_l568_c3_ac6c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node50_MUX_bit_math_h_l568_c3_ac6c_cond,
layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iftrue,
layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iffalse,
layer0_node50_MUX_bit_math_h_l568_c3_ac6c_return_output);

-- layer0_node51_MUX_bit_math_h_l579_c3_c608
layer0_node51_MUX_bit_math_h_l579_c3_c608 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node51_MUX_bit_math_h_l579_c3_c608_cond,
layer0_node51_MUX_bit_math_h_l579_c3_c608_iftrue,
layer0_node51_MUX_bit_math_h_l579_c3_c608_iffalse,
layer0_node51_MUX_bit_math_h_l579_c3_c608_return_output);

-- layer0_node52_MUX_bit_math_h_l590_c3_f975
layer0_node52_MUX_bit_math_h_l590_c3_f975 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node52_MUX_bit_math_h_l590_c3_f975_cond,
layer0_node52_MUX_bit_math_h_l590_c3_f975_iftrue,
layer0_node52_MUX_bit_math_h_l590_c3_f975_iffalse,
layer0_node52_MUX_bit_math_h_l590_c3_f975_return_output);

-- layer0_node53_MUX_bit_math_h_l601_c3_86a8
layer0_node53_MUX_bit_math_h_l601_c3_86a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node53_MUX_bit_math_h_l601_c3_86a8_cond,
layer0_node53_MUX_bit_math_h_l601_c3_86a8_iftrue,
layer0_node53_MUX_bit_math_h_l601_c3_86a8_iffalse,
layer0_node53_MUX_bit_math_h_l601_c3_86a8_return_output);

-- layer0_node54_MUX_bit_math_h_l612_c3_21f7
layer0_node54_MUX_bit_math_h_l612_c3_21f7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node54_MUX_bit_math_h_l612_c3_21f7_cond,
layer0_node54_MUX_bit_math_h_l612_c3_21f7_iftrue,
layer0_node54_MUX_bit_math_h_l612_c3_21f7_iffalse,
layer0_node54_MUX_bit_math_h_l612_c3_21f7_return_output);

-- layer0_node55_MUX_bit_math_h_l623_c3_a654
layer0_node55_MUX_bit_math_h_l623_c3_a654 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node55_MUX_bit_math_h_l623_c3_a654_cond,
layer0_node55_MUX_bit_math_h_l623_c3_a654_iftrue,
layer0_node55_MUX_bit_math_h_l623_c3_a654_iffalse,
layer0_node55_MUX_bit_math_h_l623_c3_a654_return_output);

-- layer0_node56_MUX_bit_math_h_l634_c3_259e
layer0_node56_MUX_bit_math_h_l634_c3_259e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node56_MUX_bit_math_h_l634_c3_259e_cond,
layer0_node56_MUX_bit_math_h_l634_c3_259e_iftrue,
layer0_node56_MUX_bit_math_h_l634_c3_259e_iffalse,
layer0_node56_MUX_bit_math_h_l634_c3_259e_return_output);

-- layer0_node57_MUX_bit_math_h_l645_c3_3acf
layer0_node57_MUX_bit_math_h_l645_c3_3acf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node57_MUX_bit_math_h_l645_c3_3acf_cond,
layer0_node57_MUX_bit_math_h_l645_c3_3acf_iftrue,
layer0_node57_MUX_bit_math_h_l645_c3_3acf_iffalse,
layer0_node57_MUX_bit_math_h_l645_c3_3acf_return_output);

-- layer0_node58_MUX_bit_math_h_l656_c3_6a0d
layer0_node58_MUX_bit_math_h_l656_c3_6a0d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node58_MUX_bit_math_h_l656_c3_6a0d_cond,
layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iftrue,
layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iffalse,
layer0_node58_MUX_bit_math_h_l656_c3_6a0d_return_output);

-- layer0_node59_MUX_bit_math_h_l667_c3_060a
layer0_node59_MUX_bit_math_h_l667_c3_060a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node59_MUX_bit_math_h_l667_c3_060a_cond,
layer0_node59_MUX_bit_math_h_l667_c3_060a_iftrue,
layer0_node59_MUX_bit_math_h_l667_c3_060a_iffalse,
layer0_node59_MUX_bit_math_h_l667_c3_060a_return_output);

-- layer0_node60_MUX_bit_math_h_l678_c3_dedf
layer0_node60_MUX_bit_math_h_l678_c3_dedf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node60_MUX_bit_math_h_l678_c3_dedf_cond,
layer0_node60_MUX_bit_math_h_l678_c3_dedf_iftrue,
layer0_node60_MUX_bit_math_h_l678_c3_dedf_iffalse,
layer0_node60_MUX_bit_math_h_l678_c3_dedf_return_output);

-- layer0_node61_MUX_bit_math_h_l689_c3_26a3
layer0_node61_MUX_bit_math_h_l689_c3_26a3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node61_MUX_bit_math_h_l689_c3_26a3_cond,
layer0_node61_MUX_bit_math_h_l689_c3_26a3_iftrue,
layer0_node61_MUX_bit_math_h_l689_c3_26a3_iffalse,
layer0_node61_MUX_bit_math_h_l689_c3_26a3_return_output);

-- layer0_node62_MUX_bit_math_h_l700_c3_7046
layer0_node62_MUX_bit_math_h_l700_c3_7046 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node62_MUX_bit_math_h_l700_c3_7046_cond,
layer0_node62_MUX_bit_math_h_l700_c3_7046_iftrue,
layer0_node62_MUX_bit_math_h_l700_c3_7046_iffalse,
layer0_node62_MUX_bit_math_h_l700_c3_7046_return_output);

-- layer0_node63_MUX_bit_math_h_l711_c3_0125
layer0_node63_MUX_bit_math_h_l711_c3_0125 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer0_node63_MUX_bit_math_h_l711_c3_0125_cond,
layer0_node63_MUX_bit_math_h_l711_c3_0125_iftrue,
layer0_node63_MUX_bit_math_h_l711_c3_0125_iffalse,
layer0_node63_MUX_bit_math_h_l711_c3_0125_return_output);

-- layer1_node0_MUX_bit_math_h_l728_c3_287e
layer1_node0_MUX_bit_math_h_l728_c3_287e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l728_c3_287e_cond,
layer1_node0_MUX_bit_math_h_l728_c3_287e_iftrue,
layer1_node0_MUX_bit_math_h_l728_c3_287e_iffalse,
layer1_node0_MUX_bit_math_h_l728_c3_287e_return_output);

-- layer1_node1_MUX_bit_math_h_l739_c3_3eb3
layer1_node1_MUX_bit_math_h_l739_c3_3eb3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l739_c3_3eb3_cond,
layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iftrue,
layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iffalse,
layer1_node1_MUX_bit_math_h_l739_c3_3eb3_return_output);

-- layer1_node2_MUX_bit_math_h_l750_c3_e4a0
layer1_node2_MUX_bit_math_h_l750_c3_e4a0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l750_c3_e4a0_cond,
layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iftrue,
layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iffalse,
layer1_node2_MUX_bit_math_h_l750_c3_e4a0_return_output);

-- layer1_node3_MUX_bit_math_h_l761_c3_123f
layer1_node3_MUX_bit_math_h_l761_c3_123f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l761_c3_123f_cond,
layer1_node3_MUX_bit_math_h_l761_c3_123f_iftrue,
layer1_node3_MUX_bit_math_h_l761_c3_123f_iffalse,
layer1_node3_MUX_bit_math_h_l761_c3_123f_return_output);

-- layer1_node4_MUX_bit_math_h_l772_c3_0289
layer1_node4_MUX_bit_math_h_l772_c3_0289 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node4_MUX_bit_math_h_l772_c3_0289_cond,
layer1_node4_MUX_bit_math_h_l772_c3_0289_iftrue,
layer1_node4_MUX_bit_math_h_l772_c3_0289_iffalse,
layer1_node4_MUX_bit_math_h_l772_c3_0289_return_output);

-- layer1_node5_MUX_bit_math_h_l783_c3_58a8
layer1_node5_MUX_bit_math_h_l783_c3_58a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node5_MUX_bit_math_h_l783_c3_58a8_cond,
layer1_node5_MUX_bit_math_h_l783_c3_58a8_iftrue,
layer1_node5_MUX_bit_math_h_l783_c3_58a8_iffalse,
layer1_node5_MUX_bit_math_h_l783_c3_58a8_return_output);

-- layer1_node6_MUX_bit_math_h_l794_c3_ebf4
layer1_node6_MUX_bit_math_h_l794_c3_ebf4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node6_MUX_bit_math_h_l794_c3_ebf4_cond,
layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iftrue,
layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iffalse,
layer1_node6_MUX_bit_math_h_l794_c3_ebf4_return_output);

-- layer1_node7_MUX_bit_math_h_l805_c3_1224
layer1_node7_MUX_bit_math_h_l805_c3_1224 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node7_MUX_bit_math_h_l805_c3_1224_cond,
layer1_node7_MUX_bit_math_h_l805_c3_1224_iftrue,
layer1_node7_MUX_bit_math_h_l805_c3_1224_iffalse,
layer1_node7_MUX_bit_math_h_l805_c3_1224_return_output);

-- layer1_node8_MUX_bit_math_h_l816_c3_db42
layer1_node8_MUX_bit_math_h_l816_c3_db42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node8_MUX_bit_math_h_l816_c3_db42_cond,
layer1_node8_MUX_bit_math_h_l816_c3_db42_iftrue,
layer1_node8_MUX_bit_math_h_l816_c3_db42_iffalse,
layer1_node8_MUX_bit_math_h_l816_c3_db42_return_output);

-- layer1_node9_MUX_bit_math_h_l827_c3_8290
layer1_node9_MUX_bit_math_h_l827_c3_8290 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node9_MUX_bit_math_h_l827_c3_8290_cond,
layer1_node9_MUX_bit_math_h_l827_c3_8290_iftrue,
layer1_node9_MUX_bit_math_h_l827_c3_8290_iffalse,
layer1_node9_MUX_bit_math_h_l827_c3_8290_return_output);

-- layer1_node10_MUX_bit_math_h_l838_c3_a2e2
layer1_node10_MUX_bit_math_h_l838_c3_a2e2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node10_MUX_bit_math_h_l838_c3_a2e2_cond,
layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iftrue,
layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iffalse,
layer1_node10_MUX_bit_math_h_l838_c3_a2e2_return_output);

-- layer1_node11_MUX_bit_math_h_l849_c3_dc54
layer1_node11_MUX_bit_math_h_l849_c3_dc54 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node11_MUX_bit_math_h_l849_c3_dc54_cond,
layer1_node11_MUX_bit_math_h_l849_c3_dc54_iftrue,
layer1_node11_MUX_bit_math_h_l849_c3_dc54_iffalse,
layer1_node11_MUX_bit_math_h_l849_c3_dc54_return_output);

-- layer1_node12_MUX_bit_math_h_l860_c3_7af8
layer1_node12_MUX_bit_math_h_l860_c3_7af8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node12_MUX_bit_math_h_l860_c3_7af8_cond,
layer1_node12_MUX_bit_math_h_l860_c3_7af8_iftrue,
layer1_node12_MUX_bit_math_h_l860_c3_7af8_iffalse,
layer1_node12_MUX_bit_math_h_l860_c3_7af8_return_output);

-- layer1_node13_MUX_bit_math_h_l871_c3_d1fd
layer1_node13_MUX_bit_math_h_l871_c3_d1fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node13_MUX_bit_math_h_l871_c3_d1fd_cond,
layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iftrue,
layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iffalse,
layer1_node13_MUX_bit_math_h_l871_c3_d1fd_return_output);

-- layer1_node14_MUX_bit_math_h_l882_c3_10cf
layer1_node14_MUX_bit_math_h_l882_c3_10cf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node14_MUX_bit_math_h_l882_c3_10cf_cond,
layer1_node14_MUX_bit_math_h_l882_c3_10cf_iftrue,
layer1_node14_MUX_bit_math_h_l882_c3_10cf_iffalse,
layer1_node14_MUX_bit_math_h_l882_c3_10cf_return_output);

-- layer1_node15_MUX_bit_math_h_l893_c3_3f51
layer1_node15_MUX_bit_math_h_l893_c3_3f51 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node15_MUX_bit_math_h_l893_c3_3f51_cond,
layer1_node15_MUX_bit_math_h_l893_c3_3f51_iftrue,
layer1_node15_MUX_bit_math_h_l893_c3_3f51_iffalse,
layer1_node15_MUX_bit_math_h_l893_c3_3f51_return_output);

-- layer1_node16_MUX_bit_math_h_l904_c3_e9a5
layer1_node16_MUX_bit_math_h_l904_c3_e9a5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node16_MUX_bit_math_h_l904_c3_e9a5_cond,
layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iftrue,
layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iffalse,
layer1_node16_MUX_bit_math_h_l904_c3_e9a5_return_output);

-- layer1_node17_MUX_bit_math_h_l915_c3_4b4e
layer1_node17_MUX_bit_math_h_l915_c3_4b4e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node17_MUX_bit_math_h_l915_c3_4b4e_cond,
layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iftrue,
layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iffalse,
layer1_node17_MUX_bit_math_h_l915_c3_4b4e_return_output);

-- layer1_node18_MUX_bit_math_h_l926_c3_5844
layer1_node18_MUX_bit_math_h_l926_c3_5844 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node18_MUX_bit_math_h_l926_c3_5844_cond,
layer1_node18_MUX_bit_math_h_l926_c3_5844_iftrue,
layer1_node18_MUX_bit_math_h_l926_c3_5844_iffalse,
layer1_node18_MUX_bit_math_h_l926_c3_5844_return_output);

-- layer1_node19_MUX_bit_math_h_l937_c3_7dba
layer1_node19_MUX_bit_math_h_l937_c3_7dba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node19_MUX_bit_math_h_l937_c3_7dba_cond,
layer1_node19_MUX_bit_math_h_l937_c3_7dba_iftrue,
layer1_node19_MUX_bit_math_h_l937_c3_7dba_iffalse,
layer1_node19_MUX_bit_math_h_l937_c3_7dba_return_output);

-- layer1_node20_MUX_bit_math_h_l948_c3_2725
layer1_node20_MUX_bit_math_h_l948_c3_2725 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node20_MUX_bit_math_h_l948_c3_2725_cond,
layer1_node20_MUX_bit_math_h_l948_c3_2725_iftrue,
layer1_node20_MUX_bit_math_h_l948_c3_2725_iffalse,
layer1_node20_MUX_bit_math_h_l948_c3_2725_return_output);

-- layer1_node21_MUX_bit_math_h_l959_c3_8499
layer1_node21_MUX_bit_math_h_l959_c3_8499 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node21_MUX_bit_math_h_l959_c3_8499_cond,
layer1_node21_MUX_bit_math_h_l959_c3_8499_iftrue,
layer1_node21_MUX_bit_math_h_l959_c3_8499_iffalse,
layer1_node21_MUX_bit_math_h_l959_c3_8499_return_output);

-- layer1_node22_MUX_bit_math_h_l970_c3_65bd
layer1_node22_MUX_bit_math_h_l970_c3_65bd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node22_MUX_bit_math_h_l970_c3_65bd_cond,
layer1_node22_MUX_bit_math_h_l970_c3_65bd_iftrue,
layer1_node22_MUX_bit_math_h_l970_c3_65bd_iffalse,
layer1_node22_MUX_bit_math_h_l970_c3_65bd_return_output);

-- layer1_node23_MUX_bit_math_h_l981_c3_3335
layer1_node23_MUX_bit_math_h_l981_c3_3335 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node23_MUX_bit_math_h_l981_c3_3335_cond,
layer1_node23_MUX_bit_math_h_l981_c3_3335_iftrue,
layer1_node23_MUX_bit_math_h_l981_c3_3335_iffalse,
layer1_node23_MUX_bit_math_h_l981_c3_3335_return_output);

-- layer1_node24_MUX_bit_math_h_l992_c3_8ee7
layer1_node24_MUX_bit_math_h_l992_c3_8ee7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node24_MUX_bit_math_h_l992_c3_8ee7_cond,
layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iftrue,
layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iffalse,
layer1_node24_MUX_bit_math_h_l992_c3_8ee7_return_output);

-- layer1_node25_MUX_bit_math_h_l1003_c3_8e94
layer1_node25_MUX_bit_math_h_l1003_c3_8e94 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node25_MUX_bit_math_h_l1003_c3_8e94_cond,
layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iftrue,
layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iffalse,
layer1_node25_MUX_bit_math_h_l1003_c3_8e94_return_output);

-- layer1_node26_MUX_bit_math_h_l1014_c3_d8aa
layer1_node26_MUX_bit_math_h_l1014_c3_d8aa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_cond,
layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iftrue,
layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iffalse,
layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_return_output);

-- layer1_node27_MUX_bit_math_h_l1025_c3_465f
layer1_node27_MUX_bit_math_h_l1025_c3_465f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node27_MUX_bit_math_h_l1025_c3_465f_cond,
layer1_node27_MUX_bit_math_h_l1025_c3_465f_iftrue,
layer1_node27_MUX_bit_math_h_l1025_c3_465f_iffalse,
layer1_node27_MUX_bit_math_h_l1025_c3_465f_return_output);

-- layer1_node28_MUX_bit_math_h_l1036_c3_f568
layer1_node28_MUX_bit_math_h_l1036_c3_f568 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node28_MUX_bit_math_h_l1036_c3_f568_cond,
layer1_node28_MUX_bit_math_h_l1036_c3_f568_iftrue,
layer1_node28_MUX_bit_math_h_l1036_c3_f568_iffalse,
layer1_node28_MUX_bit_math_h_l1036_c3_f568_return_output);

-- layer1_node29_MUX_bit_math_h_l1047_c3_8f77
layer1_node29_MUX_bit_math_h_l1047_c3_8f77 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node29_MUX_bit_math_h_l1047_c3_8f77_cond,
layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iftrue,
layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iffalse,
layer1_node29_MUX_bit_math_h_l1047_c3_8f77_return_output);

-- layer1_node30_MUX_bit_math_h_l1058_c3_d4dc
layer1_node30_MUX_bit_math_h_l1058_c3_d4dc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_cond,
layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iftrue,
layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iffalse,
layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_return_output);

-- layer1_node31_MUX_bit_math_h_l1069_c3_6881
layer1_node31_MUX_bit_math_h_l1069_c3_6881 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer1_node31_MUX_bit_math_h_l1069_c3_6881_cond,
layer1_node31_MUX_bit_math_h_l1069_c3_6881_iftrue,
layer1_node31_MUX_bit_math_h_l1069_c3_6881_iffalse,
layer1_node31_MUX_bit_math_h_l1069_c3_6881_return_output);

-- layer2_node0_MUX_bit_math_h_l1086_c3_f1d8
layer2_node0_MUX_bit_math_h_l1086_c3_f1d8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_cond,
layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iftrue,
layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iffalse,
layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_return_output);

-- layer2_node1_MUX_bit_math_h_l1097_c3_1a30
layer2_node1_MUX_bit_math_h_l1097_c3_1a30 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l1097_c3_1a30_cond,
layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iftrue,
layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iffalse,
layer2_node1_MUX_bit_math_h_l1097_c3_1a30_return_output);

-- layer2_node2_MUX_bit_math_h_l1108_c3_0b56
layer2_node2_MUX_bit_math_h_l1108_c3_0b56 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node2_MUX_bit_math_h_l1108_c3_0b56_cond,
layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iftrue,
layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iffalse,
layer2_node2_MUX_bit_math_h_l1108_c3_0b56_return_output);

-- layer2_node3_MUX_bit_math_h_l1119_c3_7df6
layer2_node3_MUX_bit_math_h_l1119_c3_7df6 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node3_MUX_bit_math_h_l1119_c3_7df6_cond,
layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iftrue,
layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iffalse,
layer2_node3_MUX_bit_math_h_l1119_c3_7df6_return_output);

-- layer2_node4_MUX_bit_math_h_l1130_c3_7e5b
layer2_node4_MUX_bit_math_h_l1130_c3_7e5b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_cond,
layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iftrue,
layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iffalse,
layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_return_output);

-- layer2_node5_MUX_bit_math_h_l1141_c3_25de
layer2_node5_MUX_bit_math_h_l1141_c3_25de : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node5_MUX_bit_math_h_l1141_c3_25de_cond,
layer2_node5_MUX_bit_math_h_l1141_c3_25de_iftrue,
layer2_node5_MUX_bit_math_h_l1141_c3_25de_iffalse,
layer2_node5_MUX_bit_math_h_l1141_c3_25de_return_output);

-- layer2_node6_MUX_bit_math_h_l1152_c3_be62
layer2_node6_MUX_bit_math_h_l1152_c3_be62 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node6_MUX_bit_math_h_l1152_c3_be62_cond,
layer2_node6_MUX_bit_math_h_l1152_c3_be62_iftrue,
layer2_node6_MUX_bit_math_h_l1152_c3_be62_iffalse,
layer2_node6_MUX_bit_math_h_l1152_c3_be62_return_output);

-- layer2_node7_MUX_bit_math_h_l1163_c3_9403
layer2_node7_MUX_bit_math_h_l1163_c3_9403 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node7_MUX_bit_math_h_l1163_c3_9403_cond,
layer2_node7_MUX_bit_math_h_l1163_c3_9403_iftrue,
layer2_node7_MUX_bit_math_h_l1163_c3_9403_iffalse,
layer2_node7_MUX_bit_math_h_l1163_c3_9403_return_output);

-- layer2_node8_MUX_bit_math_h_l1174_c3_918c
layer2_node8_MUX_bit_math_h_l1174_c3_918c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node8_MUX_bit_math_h_l1174_c3_918c_cond,
layer2_node8_MUX_bit_math_h_l1174_c3_918c_iftrue,
layer2_node8_MUX_bit_math_h_l1174_c3_918c_iffalse,
layer2_node8_MUX_bit_math_h_l1174_c3_918c_return_output);

-- layer2_node9_MUX_bit_math_h_l1185_c3_9e4b
layer2_node9_MUX_bit_math_h_l1185_c3_9e4b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_cond,
layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iftrue,
layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iffalse,
layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_return_output);

-- layer2_node10_MUX_bit_math_h_l1196_c3_3974
layer2_node10_MUX_bit_math_h_l1196_c3_3974 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node10_MUX_bit_math_h_l1196_c3_3974_cond,
layer2_node10_MUX_bit_math_h_l1196_c3_3974_iftrue,
layer2_node10_MUX_bit_math_h_l1196_c3_3974_iffalse,
layer2_node10_MUX_bit_math_h_l1196_c3_3974_return_output);

-- layer2_node11_MUX_bit_math_h_l1207_c3_80d7
layer2_node11_MUX_bit_math_h_l1207_c3_80d7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node11_MUX_bit_math_h_l1207_c3_80d7_cond,
layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iftrue,
layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iffalse,
layer2_node11_MUX_bit_math_h_l1207_c3_80d7_return_output);

-- layer2_node12_MUX_bit_math_h_l1218_c3_fc60
layer2_node12_MUX_bit_math_h_l1218_c3_fc60 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node12_MUX_bit_math_h_l1218_c3_fc60_cond,
layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iftrue,
layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iffalse,
layer2_node12_MUX_bit_math_h_l1218_c3_fc60_return_output);

-- layer2_node13_MUX_bit_math_h_l1229_c3_6c25
layer2_node13_MUX_bit_math_h_l1229_c3_6c25 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node13_MUX_bit_math_h_l1229_c3_6c25_cond,
layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iftrue,
layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iffalse,
layer2_node13_MUX_bit_math_h_l1229_c3_6c25_return_output);

-- layer2_node14_MUX_bit_math_h_l1240_c3_75b9
layer2_node14_MUX_bit_math_h_l1240_c3_75b9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node14_MUX_bit_math_h_l1240_c3_75b9_cond,
layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iftrue,
layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iffalse,
layer2_node14_MUX_bit_math_h_l1240_c3_75b9_return_output);

-- layer2_node15_MUX_bit_math_h_l1251_c3_ecd2
layer2_node15_MUX_bit_math_h_l1251_c3_ecd2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_cond,
layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iftrue,
layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iffalse,
layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_return_output);

-- layer3_node0_MUX_bit_math_h_l1268_c3_324b
layer3_node0_MUX_bit_math_h_l1268_c3_324b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l1268_c3_324b_cond,
layer3_node0_MUX_bit_math_h_l1268_c3_324b_iftrue,
layer3_node0_MUX_bit_math_h_l1268_c3_324b_iffalse,
layer3_node0_MUX_bit_math_h_l1268_c3_324b_return_output);

-- layer3_node1_MUX_bit_math_h_l1279_c3_eea1
layer3_node1_MUX_bit_math_h_l1279_c3_eea1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node1_MUX_bit_math_h_l1279_c3_eea1_cond,
layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iftrue,
layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iffalse,
layer3_node1_MUX_bit_math_h_l1279_c3_eea1_return_output);

-- layer3_node2_MUX_bit_math_h_l1290_c3_c56d
layer3_node2_MUX_bit_math_h_l1290_c3_c56d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node2_MUX_bit_math_h_l1290_c3_c56d_cond,
layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iftrue,
layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iffalse,
layer3_node2_MUX_bit_math_h_l1290_c3_c56d_return_output);

-- layer3_node3_MUX_bit_math_h_l1301_c3_98b1
layer3_node3_MUX_bit_math_h_l1301_c3_98b1 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node3_MUX_bit_math_h_l1301_c3_98b1_cond,
layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iftrue,
layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iffalse,
layer3_node3_MUX_bit_math_h_l1301_c3_98b1_return_output);

-- layer3_node4_MUX_bit_math_h_l1312_c3_4b99
layer3_node4_MUX_bit_math_h_l1312_c3_4b99 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node4_MUX_bit_math_h_l1312_c3_4b99_cond,
layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iftrue,
layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iffalse,
layer3_node4_MUX_bit_math_h_l1312_c3_4b99_return_output);

-- layer3_node5_MUX_bit_math_h_l1323_c3_75a2
layer3_node5_MUX_bit_math_h_l1323_c3_75a2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node5_MUX_bit_math_h_l1323_c3_75a2_cond,
layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iftrue,
layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iffalse,
layer3_node5_MUX_bit_math_h_l1323_c3_75a2_return_output);

-- layer3_node6_MUX_bit_math_h_l1334_c3_483e
layer3_node6_MUX_bit_math_h_l1334_c3_483e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node6_MUX_bit_math_h_l1334_c3_483e_cond,
layer3_node6_MUX_bit_math_h_l1334_c3_483e_iftrue,
layer3_node6_MUX_bit_math_h_l1334_c3_483e_iffalse,
layer3_node6_MUX_bit_math_h_l1334_c3_483e_return_output);

-- layer3_node7_MUX_bit_math_h_l1345_c3_7c85
layer3_node7_MUX_bit_math_h_l1345_c3_7c85 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer3_node7_MUX_bit_math_h_l1345_c3_7c85_cond,
layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iftrue,
layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iffalse,
layer3_node7_MUX_bit_math_h_l1345_c3_7c85_return_output);

-- layer4_node0_MUX_bit_math_h_l1362_c3_bbba
layer4_node0_MUX_bit_math_h_l1362_c3_bbba : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node0_MUX_bit_math_h_l1362_c3_bbba_cond,
layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iftrue,
layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iffalse,
layer4_node0_MUX_bit_math_h_l1362_c3_bbba_return_output);

-- layer4_node1_MUX_bit_math_h_l1373_c3_31df
layer4_node1_MUX_bit_math_h_l1373_c3_31df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node1_MUX_bit_math_h_l1373_c3_31df_cond,
layer4_node1_MUX_bit_math_h_l1373_c3_31df_iftrue,
layer4_node1_MUX_bit_math_h_l1373_c3_31df_iffalse,
layer4_node1_MUX_bit_math_h_l1373_c3_31df_return_output);

-- layer4_node2_MUX_bit_math_h_l1384_c3_d801
layer4_node2_MUX_bit_math_h_l1384_c3_d801 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node2_MUX_bit_math_h_l1384_c3_d801_cond,
layer4_node2_MUX_bit_math_h_l1384_c3_d801_iftrue,
layer4_node2_MUX_bit_math_h_l1384_c3_d801_iffalse,
layer4_node2_MUX_bit_math_h_l1384_c3_d801_return_output);

-- layer4_node3_MUX_bit_math_h_l1395_c3_fa88
layer4_node3_MUX_bit_math_h_l1395_c3_fa88 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer4_node3_MUX_bit_math_h_l1395_c3_fa88_cond,
layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iftrue,
layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iffalse,
layer4_node3_MUX_bit_math_h_l1395_c3_fa88_return_output);

-- layer5_node0_MUX_bit_math_h_l1412_c3_ee13
layer5_node0_MUX_bit_math_h_l1412_c3_ee13 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node0_MUX_bit_math_h_l1412_c3_ee13_cond,
layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iftrue,
layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iffalse,
layer5_node0_MUX_bit_math_h_l1412_c3_ee13_return_output);

-- layer5_node1_MUX_bit_math_h_l1423_c3_93d3
layer5_node1_MUX_bit_math_h_l1423_c3_93d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer5_node1_MUX_bit_math_h_l1423_c3_93d3_cond,
layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iftrue,
layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iffalse,
layer5_node1_MUX_bit_math_h_l1423_c3_93d3_return_output);

-- layer6_node0_MUX_bit_math_h_l1440_c3_08eb
layer6_node0_MUX_bit_math_h_l1440_c3_08eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
layer6_node0_MUX_bit_math_h_l1440_c3_08eb_cond,
layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iftrue,
layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iffalse,
layer6_node0_MUX_bit_math_h_l1440_c3_08eb_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 in16,
 in17,
 in18,
 in19,
 in20,
 in21,
 in22,
 in23,
 in24,
 in25,
 in26,
 in27,
 in28,
 in29,
 in30,
 in31,
 in32,
 in33,
 in34,
 in35,
 in36,
 in37,
 in38,
 in39,
 in40,
 in41,
 in42,
 in43,
 in44,
 in45,
 in46,
 in47,
 in48,
 in49,
 in50,
 in51,
 in52,
 in53,
 in54,
 in55,
 in56,
 in57,
 in58,
 in59,
 in60,
 in61,
 in62,
 in63,
 in64,
 in65,
 in66,
 in67,
 in68,
 in69,
 in70,
 in71,
 in72,
 in73,
 in74,
 in75,
 in76,
 in77,
 in78,
 in79,
 in80,
 in81,
 in82,
 in83,
 in84,
 in85,
 in86,
 in87,
 in88,
 in89,
 in90,
 in91,
 in92,
 in93,
 in94,
 in95,
 in96,
 in97,
 in98,
 in99,
 in100,
 in101,
 in102,
 in103,
 in104,
 in105,
 in106,
 in107,
 in108,
 in109,
 in110,
 in111,
 in112,
 in113,
 in114,
 in115,
 in116,
 in117,
 in118,
 in119,
 in120,
 in121,
 in122,
 in123,
 in124,
 in125,
 in126,
 in127,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_85c1_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_a7d4_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_43b7_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_a274_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_2eec_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_5736_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_62aa_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_c2e4_return_output,
 layer0_node8_MUX_bit_math_h_l106_c3_22f1_return_output,
 layer0_node9_MUX_bit_math_h_l117_c3_391b_return_output,
 layer0_node10_MUX_bit_math_h_l128_c3_1e58_return_output,
 layer0_node11_MUX_bit_math_h_l139_c3_6d2d_return_output,
 layer0_node12_MUX_bit_math_h_l150_c3_40e1_return_output,
 layer0_node13_MUX_bit_math_h_l161_c3_28f7_return_output,
 layer0_node14_MUX_bit_math_h_l172_c3_e31d_return_output,
 layer0_node15_MUX_bit_math_h_l183_c3_313e_return_output,
 layer0_node16_MUX_bit_math_h_l194_c3_614a_return_output,
 layer0_node17_MUX_bit_math_h_l205_c3_ec06_return_output,
 layer0_node18_MUX_bit_math_h_l216_c3_7962_return_output,
 layer0_node19_MUX_bit_math_h_l227_c3_0da7_return_output,
 layer0_node20_MUX_bit_math_h_l238_c3_a0ec_return_output,
 layer0_node21_MUX_bit_math_h_l249_c3_a3f0_return_output,
 layer0_node22_MUX_bit_math_h_l260_c3_50aa_return_output,
 layer0_node23_MUX_bit_math_h_l271_c3_b2cd_return_output,
 layer0_node24_MUX_bit_math_h_l282_c3_0847_return_output,
 layer0_node25_MUX_bit_math_h_l293_c3_d8bb_return_output,
 layer0_node26_MUX_bit_math_h_l304_c3_809a_return_output,
 layer0_node27_MUX_bit_math_h_l315_c3_a6a8_return_output,
 layer0_node28_MUX_bit_math_h_l326_c3_b62d_return_output,
 layer0_node29_MUX_bit_math_h_l337_c3_1d84_return_output,
 layer0_node30_MUX_bit_math_h_l348_c3_27f8_return_output,
 layer0_node31_MUX_bit_math_h_l359_c3_e962_return_output,
 layer0_node32_MUX_bit_math_h_l370_c3_45be_return_output,
 layer0_node33_MUX_bit_math_h_l381_c3_2a50_return_output,
 layer0_node34_MUX_bit_math_h_l392_c3_7b48_return_output,
 layer0_node35_MUX_bit_math_h_l403_c3_37e5_return_output,
 layer0_node36_MUX_bit_math_h_l414_c3_fd1a_return_output,
 layer0_node37_MUX_bit_math_h_l425_c3_8edb_return_output,
 layer0_node38_MUX_bit_math_h_l436_c3_b87e_return_output,
 layer0_node39_MUX_bit_math_h_l447_c3_8780_return_output,
 layer0_node40_MUX_bit_math_h_l458_c3_a82d_return_output,
 layer0_node41_MUX_bit_math_h_l469_c3_f332_return_output,
 layer0_node42_MUX_bit_math_h_l480_c3_8296_return_output,
 layer0_node43_MUX_bit_math_h_l491_c3_a5e9_return_output,
 layer0_node44_MUX_bit_math_h_l502_c3_7ff6_return_output,
 layer0_node45_MUX_bit_math_h_l513_c3_1806_return_output,
 layer0_node46_MUX_bit_math_h_l524_c3_c07c_return_output,
 layer0_node47_MUX_bit_math_h_l535_c3_a2fb_return_output,
 layer0_node48_MUX_bit_math_h_l546_c3_a700_return_output,
 layer0_node49_MUX_bit_math_h_l557_c3_5e53_return_output,
 layer0_node50_MUX_bit_math_h_l568_c3_ac6c_return_output,
 layer0_node51_MUX_bit_math_h_l579_c3_c608_return_output,
 layer0_node52_MUX_bit_math_h_l590_c3_f975_return_output,
 layer0_node53_MUX_bit_math_h_l601_c3_86a8_return_output,
 layer0_node54_MUX_bit_math_h_l612_c3_21f7_return_output,
 layer0_node55_MUX_bit_math_h_l623_c3_a654_return_output,
 layer0_node56_MUX_bit_math_h_l634_c3_259e_return_output,
 layer0_node57_MUX_bit_math_h_l645_c3_3acf_return_output,
 layer0_node58_MUX_bit_math_h_l656_c3_6a0d_return_output,
 layer0_node59_MUX_bit_math_h_l667_c3_060a_return_output,
 layer0_node60_MUX_bit_math_h_l678_c3_dedf_return_output,
 layer0_node61_MUX_bit_math_h_l689_c3_26a3_return_output,
 layer0_node62_MUX_bit_math_h_l700_c3_7046_return_output,
 layer0_node63_MUX_bit_math_h_l711_c3_0125_return_output,
 layer1_node0_MUX_bit_math_h_l728_c3_287e_return_output,
 layer1_node1_MUX_bit_math_h_l739_c3_3eb3_return_output,
 layer1_node2_MUX_bit_math_h_l750_c3_e4a0_return_output,
 layer1_node3_MUX_bit_math_h_l761_c3_123f_return_output,
 layer1_node4_MUX_bit_math_h_l772_c3_0289_return_output,
 layer1_node5_MUX_bit_math_h_l783_c3_58a8_return_output,
 layer1_node6_MUX_bit_math_h_l794_c3_ebf4_return_output,
 layer1_node7_MUX_bit_math_h_l805_c3_1224_return_output,
 layer1_node8_MUX_bit_math_h_l816_c3_db42_return_output,
 layer1_node9_MUX_bit_math_h_l827_c3_8290_return_output,
 layer1_node10_MUX_bit_math_h_l838_c3_a2e2_return_output,
 layer1_node11_MUX_bit_math_h_l849_c3_dc54_return_output,
 layer1_node12_MUX_bit_math_h_l860_c3_7af8_return_output,
 layer1_node13_MUX_bit_math_h_l871_c3_d1fd_return_output,
 layer1_node14_MUX_bit_math_h_l882_c3_10cf_return_output,
 layer1_node15_MUX_bit_math_h_l893_c3_3f51_return_output,
 layer1_node16_MUX_bit_math_h_l904_c3_e9a5_return_output,
 layer1_node17_MUX_bit_math_h_l915_c3_4b4e_return_output,
 layer1_node18_MUX_bit_math_h_l926_c3_5844_return_output,
 layer1_node19_MUX_bit_math_h_l937_c3_7dba_return_output,
 layer1_node20_MUX_bit_math_h_l948_c3_2725_return_output,
 layer1_node21_MUX_bit_math_h_l959_c3_8499_return_output,
 layer1_node22_MUX_bit_math_h_l970_c3_65bd_return_output,
 layer1_node23_MUX_bit_math_h_l981_c3_3335_return_output,
 layer1_node24_MUX_bit_math_h_l992_c3_8ee7_return_output,
 layer1_node25_MUX_bit_math_h_l1003_c3_8e94_return_output,
 layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_return_output,
 layer1_node27_MUX_bit_math_h_l1025_c3_465f_return_output,
 layer1_node28_MUX_bit_math_h_l1036_c3_f568_return_output,
 layer1_node29_MUX_bit_math_h_l1047_c3_8f77_return_output,
 layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_return_output,
 layer1_node31_MUX_bit_math_h_l1069_c3_6881_return_output,
 layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_return_output,
 layer2_node1_MUX_bit_math_h_l1097_c3_1a30_return_output,
 layer2_node2_MUX_bit_math_h_l1108_c3_0b56_return_output,
 layer2_node3_MUX_bit_math_h_l1119_c3_7df6_return_output,
 layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_return_output,
 layer2_node5_MUX_bit_math_h_l1141_c3_25de_return_output,
 layer2_node6_MUX_bit_math_h_l1152_c3_be62_return_output,
 layer2_node7_MUX_bit_math_h_l1163_c3_9403_return_output,
 layer2_node8_MUX_bit_math_h_l1174_c3_918c_return_output,
 layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_return_output,
 layer2_node10_MUX_bit_math_h_l1196_c3_3974_return_output,
 layer2_node11_MUX_bit_math_h_l1207_c3_80d7_return_output,
 layer2_node12_MUX_bit_math_h_l1218_c3_fc60_return_output,
 layer2_node13_MUX_bit_math_h_l1229_c3_6c25_return_output,
 layer2_node14_MUX_bit_math_h_l1240_c3_75b9_return_output,
 layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_return_output,
 layer3_node0_MUX_bit_math_h_l1268_c3_324b_return_output,
 layer3_node1_MUX_bit_math_h_l1279_c3_eea1_return_output,
 layer3_node2_MUX_bit_math_h_l1290_c3_c56d_return_output,
 layer3_node3_MUX_bit_math_h_l1301_c3_98b1_return_output,
 layer3_node4_MUX_bit_math_h_l1312_c3_4b99_return_output,
 layer3_node5_MUX_bit_math_h_l1323_c3_75a2_return_output,
 layer3_node6_MUX_bit_math_h_l1334_c3_483e_return_output,
 layer3_node7_MUX_bit_math_h_l1345_c3_7c85_return_output,
 layer4_node0_MUX_bit_math_h_l1362_c3_bbba_return_output,
 layer4_node1_MUX_bit_math_h_l1373_c3_31df_return_output,
 layer4_node2_MUX_bit_math_h_l1384_c3_d801_return_output,
 layer4_node3_MUX_bit_math_h_l1395_c3_fa88_return_output,
 layer5_node0_MUX_bit_math_h_l1412_c3_ee13_return_output,
 layer5_node1_MUX_bit_math_h_l1423_c3_93d3_return_output,
 layer6_node0_MUX_bit_math_h_l1440_c3_08eb_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(7 downto 0);
 variable VAR_sel : unsigned(6 downto 0);
 variable VAR_in0 : unsigned(7 downto 0);
 variable VAR_in1 : unsigned(7 downto 0);
 variable VAR_in2 : unsigned(7 downto 0);
 variable VAR_in3 : unsigned(7 downto 0);
 variable VAR_in4 : unsigned(7 downto 0);
 variable VAR_in5 : unsigned(7 downto 0);
 variable VAR_in6 : unsigned(7 downto 0);
 variable VAR_in7 : unsigned(7 downto 0);
 variable VAR_in8 : unsigned(7 downto 0);
 variable VAR_in9 : unsigned(7 downto 0);
 variable VAR_in10 : unsigned(7 downto 0);
 variable VAR_in11 : unsigned(7 downto 0);
 variable VAR_in12 : unsigned(7 downto 0);
 variable VAR_in13 : unsigned(7 downto 0);
 variable VAR_in14 : unsigned(7 downto 0);
 variable VAR_in15 : unsigned(7 downto 0);
 variable VAR_in16 : unsigned(7 downto 0);
 variable VAR_in17 : unsigned(7 downto 0);
 variable VAR_in18 : unsigned(7 downto 0);
 variable VAR_in19 : unsigned(7 downto 0);
 variable VAR_in20 : unsigned(7 downto 0);
 variable VAR_in21 : unsigned(7 downto 0);
 variable VAR_in22 : unsigned(7 downto 0);
 variable VAR_in23 : unsigned(7 downto 0);
 variable VAR_in24 : unsigned(7 downto 0);
 variable VAR_in25 : unsigned(7 downto 0);
 variable VAR_in26 : unsigned(7 downto 0);
 variable VAR_in27 : unsigned(7 downto 0);
 variable VAR_in28 : unsigned(7 downto 0);
 variable VAR_in29 : unsigned(7 downto 0);
 variable VAR_in30 : unsigned(7 downto 0);
 variable VAR_in31 : unsigned(7 downto 0);
 variable VAR_in32 : unsigned(7 downto 0);
 variable VAR_in33 : unsigned(7 downto 0);
 variable VAR_in34 : unsigned(7 downto 0);
 variable VAR_in35 : unsigned(7 downto 0);
 variable VAR_in36 : unsigned(7 downto 0);
 variable VAR_in37 : unsigned(7 downto 0);
 variable VAR_in38 : unsigned(7 downto 0);
 variable VAR_in39 : unsigned(7 downto 0);
 variable VAR_in40 : unsigned(7 downto 0);
 variable VAR_in41 : unsigned(7 downto 0);
 variable VAR_in42 : unsigned(7 downto 0);
 variable VAR_in43 : unsigned(7 downto 0);
 variable VAR_in44 : unsigned(7 downto 0);
 variable VAR_in45 : unsigned(7 downto 0);
 variable VAR_in46 : unsigned(7 downto 0);
 variable VAR_in47 : unsigned(7 downto 0);
 variable VAR_in48 : unsigned(7 downto 0);
 variable VAR_in49 : unsigned(7 downto 0);
 variable VAR_in50 : unsigned(7 downto 0);
 variable VAR_in51 : unsigned(7 downto 0);
 variable VAR_in52 : unsigned(7 downto 0);
 variable VAR_in53 : unsigned(7 downto 0);
 variable VAR_in54 : unsigned(7 downto 0);
 variable VAR_in55 : unsigned(7 downto 0);
 variable VAR_in56 : unsigned(7 downto 0);
 variable VAR_in57 : unsigned(7 downto 0);
 variable VAR_in58 : unsigned(7 downto 0);
 variable VAR_in59 : unsigned(7 downto 0);
 variable VAR_in60 : unsigned(7 downto 0);
 variable VAR_in61 : unsigned(7 downto 0);
 variable VAR_in62 : unsigned(7 downto 0);
 variable VAR_in63 : unsigned(7 downto 0);
 variable VAR_in64 : unsigned(7 downto 0);
 variable VAR_in65 : unsigned(7 downto 0);
 variable VAR_in66 : unsigned(7 downto 0);
 variable VAR_in67 : unsigned(7 downto 0);
 variable VAR_in68 : unsigned(7 downto 0);
 variable VAR_in69 : unsigned(7 downto 0);
 variable VAR_in70 : unsigned(7 downto 0);
 variable VAR_in71 : unsigned(7 downto 0);
 variable VAR_in72 : unsigned(7 downto 0);
 variable VAR_in73 : unsigned(7 downto 0);
 variable VAR_in74 : unsigned(7 downto 0);
 variable VAR_in75 : unsigned(7 downto 0);
 variable VAR_in76 : unsigned(7 downto 0);
 variable VAR_in77 : unsigned(7 downto 0);
 variable VAR_in78 : unsigned(7 downto 0);
 variable VAR_in79 : unsigned(7 downto 0);
 variable VAR_in80 : unsigned(7 downto 0);
 variable VAR_in81 : unsigned(7 downto 0);
 variable VAR_in82 : unsigned(7 downto 0);
 variable VAR_in83 : unsigned(7 downto 0);
 variable VAR_in84 : unsigned(7 downto 0);
 variable VAR_in85 : unsigned(7 downto 0);
 variable VAR_in86 : unsigned(7 downto 0);
 variable VAR_in87 : unsigned(7 downto 0);
 variable VAR_in88 : unsigned(7 downto 0);
 variable VAR_in89 : unsigned(7 downto 0);
 variable VAR_in90 : unsigned(7 downto 0);
 variable VAR_in91 : unsigned(7 downto 0);
 variable VAR_in92 : unsigned(7 downto 0);
 variable VAR_in93 : unsigned(7 downto 0);
 variable VAR_in94 : unsigned(7 downto 0);
 variable VAR_in95 : unsigned(7 downto 0);
 variable VAR_in96 : unsigned(7 downto 0);
 variable VAR_in97 : unsigned(7 downto 0);
 variable VAR_in98 : unsigned(7 downto 0);
 variable VAR_in99 : unsigned(7 downto 0);
 variable VAR_in100 : unsigned(7 downto 0);
 variable VAR_in101 : unsigned(7 downto 0);
 variable VAR_in102 : unsigned(7 downto 0);
 variable VAR_in103 : unsigned(7 downto 0);
 variable VAR_in104 : unsigned(7 downto 0);
 variable VAR_in105 : unsigned(7 downto 0);
 variable VAR_in106 : unsigned(7 downto 0);
 variable VAR_in107 : unsigned(7 downto 0);
 variable VAR_in108 : unsigned(7 downto 0);
 variable VAR_in109 : unsigned(7 downto 0);
 variable VAR_in110 : unsigned(7 downto 0);
 variable VAR_in111 : unsigned(7 downto 0);
 variable VAR_in112 : unsigned(7 downto 0);
 variable VAR_in113 : unsigned(7 downto 0);
 variable VAR_in114 : unsigned(7 downto 0);
 variable VAR_in115 : unsigned(7 downto 0);
 variable VAR_in116 : unsigned(7 downto 0);
 variable VAR_in117 : unsigned(7 downto 0);
 variable VAR_in118 : unsigned(7 downto 0);
 variable VAR_in119 : unsigned(7 downto 0);
 variable VAR_in120 : unsigned(7 downto 0);
 variable VAR_in121 : unsigned(7 downto 0);
 variable VAR_in122 : unsigned(7 downto 0);
 variable VAR_in123 : unsigned(7 downto 0);
 variable VAR_in124 : unsigned(7 downto 0);
 variable VAR_in125 : unsigned(7 downto 0);
 variable VAR_in126 : unsigned(7 downto 0);
 variable VAR_in127 : unsigned(7 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_cond : unsigned(0 downto 0);
 variable VAR_layer0_node8 : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node9 : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_cond : unsigned(0 downto 0);
 variable VAR_layer0_node10 : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_cond : unsigned(0 downto 0);
 variable VAR_layer0_node11 : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node12 : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_cond : unsigned(0 downto 0);
 variable VAR_layer0_node13 : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node14 : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node15 : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node16 : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node17 : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_cond : unsigned(0 downto 0);
 variable VAR_layer0_node18 : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_cond : unsigned(0 downto 0);
 variable VAR_layer0_node19 : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node20 : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_cond : unsigned(0 downto 0);
 variable VAR_layer0_node21 : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_cond : unsigned(0 downto 0);
 variable VAR_layer0_node22 : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_cond : unsigned(0 downto 0);
 variable VAR_layer0_node23 : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_cond : unsigned(0 downto 0);
 variable VAR_layer0_node24 : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_cond : unsigned(0 downto 0);
 variable VAR_layer0_node25 : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_cond : unsigned(0 downto 0);
 variable VAR_layer0_node26 : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node27 : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node28 : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node29 : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_cond : unsigned(0 downto 0);
 variable VAR_layer0_node30 : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node31 : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_cond : unsigned(0 downto 0);
 variable VAR_layer0_node32 : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_cond : unsigned(0 downto 0);
 variable VAR_layer0_node33 : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_cond : unsigned(0 downto 0);
 variable VAR_layer0_node34 : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_cond : unsigned(0 downto 0);
 variable VAR_layer0_node35 : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_cond : unsigned(0 downto 0);
 variable VAR_layer0_node36 : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node37 : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_cond : unsigned(0 downto 0);
 variable VAR_layer0_node38 : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node39 : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_cond : unsigned(0 downto 0);
 variable VAR_layer0_node40 : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node41 : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_cond : unsigned(0 downto 0);
 variable VAR_layer0_node42 : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_cond : unsigned(0 downto 0);
 variable VAR_layer0_node43 : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_cond : unsigned(0 downto 0);
 variable VAR_layer0_node44 : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_cond : unsigned(0 downto 0);
 variable VAR_layer0_node45 : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_cond : unsigned(0 downto 0);
 variable VAR_layer0_node46 : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node47 : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_cond : unsigned(0 downto 0);
 variable VAR_layer0_node48 : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_cond : unsigned(0 downto 0);
 variable VAR_layer0_node49 : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_cond : unsigned(0 downto 0);
 variable VAR_layer0_node50 : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_cond : unsigned(0 downto 0);
 variable VAR_layer0_node51 : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_cond : unsigned(0 downto 0);
 variable VAR_layer0_node52 : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_cond : unsigned(0 downto 0);
 variable VAR_layer0_node53 : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_cond : unsigned(0 downto 0);
 variable VAR_layer0_node54 : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node55 : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_cond : unsigned(0 downto 0);
 variable VAR_layer0_node56 : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_cond : unsigned(0 downto 0);
 variable VAR_layer0_node57 : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_cond : unsigned(0 downto 0);
 variable VAR_layer0_node58 : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node59 : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node60 : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_cond : unsigned(0 downto 0);
 variable VAR_layer0_node61 : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_cond : unsigned(0 downto 0);
 variable VAR_layer0_node62 : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_cond : unsigned(0 downto 0);
 variable VAR_layer0_node63 : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_iftrue : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_iffalse : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_return_output : unsigned(7 downto 0);
 variable VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node4 : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_cond : unsigned(0 downto 0);
 variable VAR_layer1_node5 : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_cond : unsigned(0 downto 0);
 variable VAR_layer1_node6 : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_cond : unsigned(0 downto 0);
 variable VAR_layer1_node7 : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_cond : unsigned(0 downto 0);
 variable VAR_layer1_node8 : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_cond : unsigned(0 downto 0);
 variable VAR_layer1_node9 : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_cond : unsigned(0 downto 0);
 variable VAR_layer1_node10 : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_cond : unsigned(0 downto 0);
 variable VAR_layer1_node11 : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_cond : unsigned(0 downto 0);
 variable VAR_layer1_node12 : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_cond : unsigned(0 downto 0);
 variable VAR_layer1_node13 : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_cond : unsigned(0 downto 0);
 variable VAR_layer1_node14 : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_cond : unsigned(0 downto 0);
 variable VAR_layer1_node15 : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_cond : unsigned(0 downto 0);
 variable VAR_layer1_node16 : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_cond : unsigned(0 downto 0);
 variable VAR_layer1_node17 : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_cond : unsigned(0 downto 0);
 variable VAR_layer1_node18 : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_cond : unsigned(0 downto 0);
 variable VAR_layer1_node19 : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_cond : unsigned(0 downto 0);
 variable VAR_layer1_node20 : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_cond : unsigned(0 downto 0);
 variable VAR_layer1_node21 : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_cond : unsigned(0 downto 0);
 variable VAR_layer1_node22 : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_cond : unsigned(0 downto 0);
 variable VAR_layer1_node23 : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_cond : unsigned(0 downto 0);
 variable VAR_layer1_node24 : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_cond : unsigned(0 downto 0);
 variable VAR_layer1_node25 : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_cond : unsigned(0 downto 0);
 variable VAR_layer1_node26 : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_cond : unsigned(0 downto 0);
 variable VAR_layer1_node27 : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_cond : unsigned(0 downto 0);
 variable VAR_layer1_node28 : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_cond : unsigned(0 downto 0);
 variable VAR_layer1_node29 : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_cond : unsigned(0 downto 0);
 variable VAR_layer1_node30 : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_cond : unsigned(0 downto 0);
 variable VAR_layer1_node31 : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_iftrue : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_iffalse : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_return_output : unsigned(7 downto 0);
 variable VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_cond : unsigned(0 downto 0);
 variable VAR_layer2_node2 : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_cond : unsigned(0 downto 0);
 variable VAR_layer2_node3 : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_cond : unsigned(0 downto 0);
 variable VAR_layer2_node4 : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_cond : unsigned(0 downto 0);
 variable VAR_layer2_node5 : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_cond : unsigned(0 downto 0);
 variable VAR_layer2_node6 : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_cond : unsigned(0 downto 0);
 variable VAR_layer2_node7 : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_cond : unsigned(0 downto 0);
 variable VAR_layer2_node8 : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_cond : unsigned(0 downto 0);
 variable VAR_layer2_node9 : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_cond : unsigned(0 downto 0);
 variable VAR_layer2_node10 : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_cond : unsigned(0 downto 0);
 variable VAR_layer2_node11 : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_cond : unsigned(0 downto 0);
 variable VAR_layer2_node12 : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_cond : unsigned(0 downto 0);
 variable VAR_layer2_node13 : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_cond : unsigned(0 downto 0);
 variable VAR_layer2_node14 : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_cond : unsigned(0 downto 0);
 variable VAR_layer2_node15 : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iftrue : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iffalse : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_return_output : unsigned(7 downto 0);
 variable VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_cond : unsigned(0 downto 0);
 variable VAR_layer3_node1 : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_cond : unsigned(0 downto 0);
 variable VAR_layer3_node2 : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_cond : unsigned(0 downto 0);
 variable VAR_layer3_node3 : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_cond : unsigned(0 downto 0);
 variable VAR_layer3_node4 : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_cond : unsigned(0 downto 0);
 variable VAR_layer3_node5 : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_cond : unsigned(0 downto 0);
 variable VAR_layer3_node6 : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_cond : unsigned(0 downto 0);
 variable VAR_layer3_node7 : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iftrue : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iffalse : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_return_output : unsigned(7 downto 0);
 variable VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_cond : unsigned(0 downto 0);
 variable VAR_sel4 : unsigned(0 downto 0);
 variable VAR_uint7_4_4_bit_math_h_l1358_c10_6da6_return_output : unsigned(0 downto 0);
 variable VAR_layer4_node0 : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_cond : unsigned(0 downto 0);
 variable VAR_layer4_node1 : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_cond : unsigned(0 downto 0);
 variable VAR_layer4_node2 : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_cond : unsigned(0 downto 0);
 variable VAR_layer4_node3 : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iftrue : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iffalse : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_return_output : unsigned(7 downto 0);
 variable VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_cond : unsigned(0 downto 0);
 variable VAR_sel5 : unsigned(0 downto 0);
 variable VAR_uint7_5_5_bit_math_h_l1408_c10_7a52_return_output : unsigned(0 downto 0);
 variable VAR_layer5_node0 : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_cond : unsigned(0 downto 0);
 variable VAR_layer5_node1 : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iftrue : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iffalse : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_return_output : unsigned(7 downto 0);
 variable VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_cond : unsigned(0 downto 0);
 variable VAR_sel6 : unsigned(0 downto 0);
 variable VAR_uint7_6_6_bit_math_h_l1436_c10_d6aa_return_output : unsigned(0 downto 0);
 variable VAR_layer6_node0 : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iftrue : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iffalse : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_return_output : unsigned(7 downto 0);
 variable VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;
     VAR_in16 := in16;
     VAR_in17 := in17;
     VAR_in18 := in18;
     VAR_in19 := in19;
     VAR_in20 := in20;
     VAR_in21 := in21;
     VAR_in22 := in22;
     VAR_in23 := in23;
     VAR_in24 := in24;
     VAR_in25 := in25;
     VAR_in26 := in26;
     VAR_in27 := in27;
     VAR_in28 := in28;
     VAR_in29 := in29;
     VAR_in30 := in30;
     VAR_in31 := in31;
     VAR_in32 := in32;
     VAR_in33 := in33;
     VAR_in34 := in34;
     VAR_in35 := in35;
     VAR_in36 := in36;
     VAR_in37 := in37;
     VAR_in38 := in38;
     VAR_in39 := in39;
     VAR_in40 := in40;
     VAR_in41 := in41;
     VAR_in42 := in42;
     VAR_in43 := in43;
     VAR_in44 := in44;
     VAR_in45 := in45;
     VAR_in46 := in46;
     VAR_in47 := in47;
     VAR_in48 := in48;
     VAR_in49 := in49;
     VAR_in50 := in50;
     VAR_in51 := in51;
     VAR_in52 := in52;
     VAR_in53 := in53;
     VAR_in54 := in54;
     VAR_in55 := in55;
     VAR_in56 := in56;
     VAR_in57 := in57;
     VAR_in58 := in58;
     VAR_in59 := in59;
     VAR_in60 := in60;
     VAR_in61 := in61;
     VAR_in62 := in62;
     VAR_in63 := in63;
     VAR_in64 := in64;
     VAR_in65 := in65;
     VAR_in66 := in66;
     VAR_in67 := in67;
     VAR_in68 := in68;
     VAR_in69 := in69;
     VAR_in70 := in70;
     VAR_in71 := in71;
     VAR_in72 := in72;
     VAR_in73 := in73;
     VAR_in74 := in74;
     VAR_in75 := in75;
     VAR_in76 := in76;
     VAR_in77 := in77;
     VAR_in78 := in78;
     VAR_in79 := in79;
     VAR_in80 := in80;
     VAR_in81 := in81;
     VAR_in82 := in82;
     VAR_in83 := in83;
     VAR_in84 := in84;
     VAR_in85 := in85;
     VAR_in86 := in86;
     VAR_in87 := in87;
     VAR_in88 := in88;
     VAR_in89 := in89;
     VAR_in90 := in90;
     VAR_in91 := in91;
     VAR_in92 := in92;
     VAR_in93 := in93;
     VAR_in94 := in94;
     VAR_in95 := in95;
     VAR_in96 := in96;
     VAR_in97 := in97;
     VAR_in98 := in98;
     VAR_in99 := in99;
     VAR_in100 := in100;
     VAR_in101 := in101;
     VAR_in102 := in102;
     VAR_in103 := in103;
     VAR_in104 := in104;
     VAR_in105 := in105;
     VAR_in106 := in106;
     VAR_in107 := in107;
     VAR_in108 := in108;
     VAR_in109 := in109;
     VAR_in110 := in110;
     VAR_in111 := in111;
     VAR_in112 := in112;
     VAR_in113 := in113;
     VAR_in114 := in114;
     VAR_in115 := in115;
     VAR_in116 := in116;
     VAR_in117 := in117;
     VAR_in118 := in118;
     VAR_in119 := in119;
     VAR_in120 := in120;
     VAR_in121 := in121;
     VAR_in122 := in122;
     VAR_in123 := in123;
     VAR_in124 := in124;
     VAR_in125 := in125;
     VAR_in126 := in126;
     VAR_in127 := in127;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_iffalse := VAR_in10;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iffalse := VAR_in100;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iftrue := VAR_in101;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_iffalse := VAR_in102;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_iftrue := VAR_in103;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_iffalse := VAR_in104;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_iftrue := VAR_in105;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_iffalse := VAR_in106;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_iftrue := VAR_in107;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_iffalse := VAR_in108;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_iftrue := VAR_in109;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_iftrue := VAR_in11;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_iffalse := VAR_in110;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_iftrue := VAR_in111;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_iffalse := VAR_in112;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_iftrue := VAR_in113;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_iffalse := VAR_in114;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_iftrue := VAR_in115;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iffalse := VAR_in116;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iftrue := VAR_in117;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_iffalse := VAR_in118;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_iftrue := VAR_in119;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_iffalse := VAR_in12;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_iffalse := VAR_in120;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_iftrue := VAR_in121;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_iffalse := VAR_in122;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_iftrue := VAR_in123;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_iffalse := VAR_in124;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_iftrue := VAR_in125;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_iffalse := VAR_in126;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_iftrue := VAR_in127;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iftrue := VAR_in15;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_iffalse := VAR_in16;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_iftrue := VAR_in17;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_iffalse := VAR_in18;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_iftrue := VAR_in19;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iffalse := VAR_in2;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_iffalse := VAR_in20;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_iftrue := VAR_in21;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iffalse := VAR_in22;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iftrue := VAR_in23;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_iffalse := VAR_in24;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_iftrue := VAR_in25;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_iffalse := VAR_in26;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_iftrue := VAR_in27;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_iffalse := VAR_in28;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_iftrue := VAR_in29;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iftrue := VAR_in3;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_iffalse := VAR_in30;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_iftrue := VAR_in31;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_iffalse := VAR_in32;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_iftrue := VAR_in33;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_iffalse := VAR_in34;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_iftrue := VAR_in35;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_iffalse := VAR_in36;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_iftrue := VAR_in37;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_iffalse := VAR_in38;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_iftrue := VAR_in39;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_iffalse := VAR_in4;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iffalse := VAR_in40;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iftrue := VAR_in41;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iffalse := VAR_in42;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iftrue := VAR_in43;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_iffalse := VAR_in44;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_iftrue := VAR_in45;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iffalse := VAR_in46;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iftrue := VAR_in47;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_iffalse := VAR_in48;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_iftrue := VAR_in49;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_iftrue := VAR_in5;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iffalse := VAR_in50;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iftrue := VAR_in51;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_iffalse := VAR_in52;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_iftrue := VAR_in53;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iffalse := VAR_in54;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iftrue := VAR_in55;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_iffalse := VAR_in56;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_iftrue := VAR_in57;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_iffalse := VAR_in58;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_iftrue := VAR_in59;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_iffalse := VAR_in6;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_iffalse := VAR_in60;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_iftrue := VAR_in61;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_iffalse := VAR_in62;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_iftrue := VAR_in63;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_iffalse := VAR_in64;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_iftrue := VAR_in65;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_iffalse := VAR_in66;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_iftrue := VAR_in67;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_iffalse := VAR_in68;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_iftrue := VAR_in69;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_iftrue := VAR_in7;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_iffalse := VAR_in70;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_iftrue := VAR_in71;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iffalse := VAR_in72;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iftrue := VAR_in73;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_iffalse := VAR_in74;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_iftrue := VAR_in75;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_iffalse := VAR_in76;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_iftrue := VAR_in77;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_iffalse := VAR_in78;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_iftrue := VAR_in79;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_iffalse := VAR_in8;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_iffalse := VAR_in80;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_iftrue := VAR_in81;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_iffalse := VAR_in82;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_iftrue := VAR_in83;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_iffalse := VAR_in84;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_iftrue := VAR_in85;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iffalse := VAR_in86;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iftrue := VAR_in87;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iffalse := VAR_in88;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iftrue := VAR_in89;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_iftrue := VAR_in9;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_iffalse := VAR_in90;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_iftrue := VAR_in91;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_iffalse := VAR_in92;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_iftrue := VAR_in93;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iffalse := VAR_in94;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iftrue := VAR_in95;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_iffalse := VAR_in96;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_iftrue := VAR_in97;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_iffalse := VAR_in98;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_iftrue := VAR_in99;
     -- uint7_1_1[bit_math_h_l724_c10_d41a] LATENCY=0
     VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output := uint7_1_1(
     VAR_sel);

     -- uint7_4_4[bit_math_h_l1358_c10_6da6] LATENCY=0
     VAR_uint7_4_4_bit_math_h_l1358_c10_6da6_return_output := uint7_4_4(
     VAR_sel);

     -- uint7_2_2[bit_math_h_l1082_c10_bd43] LATENCY=0
     VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output := uint7_2_2(
     VAR_sel);

     -- uint7_3_3[bit_math_h_l1264_c10_b672] LATENCY=0
     VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output := uint7_3_3(
     VAR_sel);

     -- uint7_6_6[bit_math_h_l1436_c10_d6aa] LATENCY=0
     VAR_uint7_6_6_bit_math_h_l1436_c10_d6aa_return_output := uint7_6_6(
     VAR_sel);

     -- uint7_0_0[bit_math_h_l14_c10_d67b] LATENCY=0
     VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output := uint7_0_0(
     VAR_sel);

     -- uint7_5_5[bit_math_h_l1408_c10_7a52] LATENCY=0
     VAR_uint7_5_5_bit_math_h_l1408_c10_7a52_return_output := uint7_5_5(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_cond := VAR_uint7_0_0_bit_math_h_l14_c10_d67b_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_cond := VAR_uint7_1_1_bit_math_h_l724_c10_d41a_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_cond := VAR_uint7_2_2_bit_math_h_l1082_c10_bd43_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_cond := VAR_uint7_3_3_bit_math_h_l1264_c10_b672_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_6da6_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_6da6_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_6da6_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_cond := VAR_uint7_4_4_bit_math_h_l1358_c10_6da6_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_7a52_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_cond := VAR_uint7_5_5_bit_math_h_l1408_c10_7a52_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_cond := VAR_uint7_6_6_bit_math_h_l1436_c10_d6aa_return_output;
     -- layer0_node1_MUX[bit_math_h_l29_c3_a7d4] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_a7d4_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_return_output := layer0_node1_MUX_bit_math_h_l29_c3_a7d4_return_output;

     -- layer0_node10_MUX[bit_math_h_l128_c3_1e58] LATENCY=0
     -- Inputs
     layer0_node10_MUX_bit_math_h_l128_c3_1e58_cond <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_cond;
     layer0_node10_MUX_bit_math_h_l128_c3_1e58_iftrue <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_iftrue;
     layer0_node10_MUX_bit_math_h_l128_c3_1e58_iffalse <= VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_iffalse;
     -- Outputs
     VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_return_output := layer0_node10_MUX_bit_math_h_l128_c3_1e58_return_output;

     -- layer0_node11_MUX[bit_math_h_l139_c3_6d2d] LATENCY=0
     -- Inputs
     layer0_node11_MUX_bit_math_h_l139_c3_6d2d_cond <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_cond;
     layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iftrue <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iftrue;
     layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iffalse <= VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_iffalse;
     -- Outputs
     VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_return_output := layer0_node11_MUX_bit_math_h_l139_c3_6d2d_return_output;

     -- layer0_node13_MUX[bit_math_h_l161_c3_28f7] LATENCY=0
     -- Inputs
     layer0_node13_MUX_bit_math_h_l161_c3_28f7_cond <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_cond;
     layer0_node13_MUX_bit_math_h_l161_c3_28f7_iftrue <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_iftrue;
     layer0_node13_MUX_bit_math_h_l161_c3_28f7_iffalse <= VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_iffalse;
     -- Outputs
     VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_return_output := layer0_node13_MUX_bit_math_h_l161_c3_28f7_return_output;

     -- layer0_node41_MUX[bit_math_h_l469_c3_f332] LATENCY=0
     -- Inputs
     layer0_node41_MUX_bit_math_h_l469_c3_f332_cond <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_cond;
     layer0_node41_MUX_bit_math_h_l469_c3_f332_iftrue <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_iftrue;
     layer0_node41_MUX_bit_math_h_l469_c3_f332_iffalse <= VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_iffalse;
     -- Outputs
     VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_return_output := layer0_node41_MUX_bit_math_h_l469_c3_f332_return_output;

     -- layer0_node36_MUX[bit_math_h_l414_c3_fd1a] LATENCY=0
     -- Inputs
     layer0_node36_MUX_bit_math_h_l414_c3_fd1a_cond <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_cond;
     layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iftrue <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iftrue;
     layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iffalse <= VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_iffalse;
     -- Outputs
     VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_return_output := layer0_node36_MUX_bit_math_h_l414_c3_fd1a_return_output;

     -- layer0_node61_MUX[bit_math_h_l689_c3_26a3] LATENCY=0
     -- Inputs
     layer0_node61_MUX_bit_math_h_l689_c3_26a3_cond <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_cond;
     layer0_node61_MUX_bit_math_h_l689_c3_26a3_iftrue <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_iftrue;
     layer0_node61_MUX_bit_math_h_l689_c3_26a3_iffalse <= VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_iffalse;
     -- Outputs
     VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_return_output := layer0_node61_MUX_bit_math_h_l689_c3_26a3_return_output;

     -- layer0_node48_MUX[bit_math_h_l546_c3_a700] LATENCY=0
     -- Inputs
     layer0_node48_MUX_bit_math_h_l546_c3_a700_cond <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_cond;
     layer0_node48_MUX_bit_math_h_l546_c3_a700_iftrue <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_iftrue;
     layer0_node48_MUX_bit_math_h_l546_c3_a700_iffalse <= VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_iffalse;
     -- Outputs
     VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_return_output := layer0_node48_MUX_bit_math_h_l546_c3_a700_return_output;

     -- layer0_node63_MUX[bit_math_h_l711_c3_0125] LATENCY=0
     -- Inputs
     layer0_node63_MUX_bit_math_h_l711_c3_0125_cond <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_cond;
     layer0_node63_MUX_bit_math_h_l711_c3_0125_iftrue <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_iftrue;
     layer0_node63_MUX_bit_math_h_l711_c3_0125_iffalse <= VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_iffalse;
     -- Outputs
     VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_return_output := layer0_node63_MUX_bit_math_h_l711_c3_0125_return_output;

     -- layer0_node39_MUX[bit_math_h_l447_c3_8780] LATENCY=0
     -- Inputs
     layer0_node39_MUX_bit_math_h_l447_c3_8780_cond <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_cond;
     layer0_node39_MUX_bit_math_h_l447_c3_8780_iftrue <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_iftrue;
     layer0_node39_MUX_bit_math_h_l447_c3_8780_iffalse <= VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_iffalse;
     -- Outputs
     VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_return_output := layer0_node39_MUX_bit_math_h_l447_c3_8780_return_output;

     -- layer0_node42_MUX[bit_math_h_l480_c3_8296] LATENCY=0
     -- Inputs
     layer0_node42_MUX_bit_math_h_l480_c3_8296_cond <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_cond;
     layer0_node42_MUX_bit_math_h_l480_c3_8296_iftrue <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_iftrue;
     layer0_node42_MUX_bit_math_h_l480_c3_8296_iffalse <= VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_iffalse;
     -- Outputs
     VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_return_output := layer0_node42_MUX_bit_math_h_l480_c3_8296_return_output;

     -- layer0_node58_MUX[bit_math_h_l656_c3_6a0d] LATENCY=0
     -- Inputs
     layer0_node58_MUX_bit_math_h_l656_c3_6a0d_cond <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_cond;
     layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iftrue <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iftrue;
     layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iffalse <= VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_iffalse;
     -- Outputs
     VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_return_output := layer0_node58_MUX_bit_math_h_l656_c3_6a0d_return_output;

     -- layer0_node21_MUX[bit_math_h_l249_c3_a3f0] LATENCY=0
     -- Inputs
     layer0_node21_MUX_bit_math_h_l249_c3_a3f0_cond <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_cond;
     layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iftrue <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iftrue;
     layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iffalse <= VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_iffalse;
     -- Outputs
     VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_return_output := layer0_node21_MUX_bit_math_h_l249_c3_a3f0_return_output;

     -- layer0_node57_MUX[bit_math_h_l645_c3_3acf] LATENCY=0
     -- Inputs
     layer0_node57_MUX_bit_math_h_l645_c3_3acf_cond <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_cond;
     layer0_node57_MUX_bit_math_h_l645_c3_3acf_iftrue <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_iftrue;
     layer0_node57_MUX_bit_math_h_l645_c3_3acf_iffalse <= VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_iffalse;
     -- Outputs
     VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_return_output := layer0_node57_MUX_bit_math_h_l645_c3_3acf_return_output;

     -- layer0_node12_MUX[bit_math_h_l150_c3_40e1] LATENCY=0
     -- Inputs
     layer0_node12_MUX_bit_math_h_l150_c3_40e1_cond <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_cond;
     layer0_node12_MUX_bit_math_h_l150_c3_40e1_iftrue <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_iftrue;
     layer0_node12_MUX_bit_math_h_l150_c3_40e1_iffalse <= VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_iffalse;
     -- Outputs
     VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_return_output := layer0_node12_MUX_bit_math_h_l150_c3_40e1_return_output;

     -- layer0_node28_MUX[bit_math_h_l326_c3_b62d] LATENCY=0
     -- Inputs
     layer0_node28_MUX_bit_math_h_l326_c3_b62d_cond <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_cond;
     layer0_node28_MUX_bit_math_h_l326_c3_b62d_iftrue <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_iftrue;
     layer0_node28_MUX_bit_math_h_l326_c3_b62d_iffalse <= VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_iffalse;
     -- Outputs
     VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_return_output := layer0_node28_MUX_bit_math_h_l326_c3_b62d_return_output;

     -- layer0_node16_MUX[bit_math_h_l194_c3_614a] LATENCY=0
     -- Inputs
     layer0_node16_MUX_bit_math_h_l194_c3_614a_cond <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_cond;
     layer0_node16_MUX_bit_math_h_l194_c3_614a_iftrue <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_iftrue;
     layer0_node16_MUX_bit_math_h_l194_c3_614a_iffalse <= VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_iffalse;
     -- Outputs
     VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_return_output := layer0_node16_MUX_bit_math_h_l194_c3_614a_return_output;

     -- layer0_node37_MUX[bit_math_h_l425_c3_8edb] LATENCY=0
     -- Inputs
     layer0_node37_MUX_bit_math_h_l425_c3_8edb_cond <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_cond;
     layer0_node37_MUX_bit_math_h_l425_c3_8edb_iftrue <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_iftrue;
     layer0_node37_MUX_bit_math_h_l425_c3_8edb_iffalse <= VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_iffalse;
     -- Outputs
     VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_return_output := layer0_node37_MUX_bit_math_h_l425_c3_8edb_return_output;

     -- layer0_node51_MUX[bit_math_h_l579_c3_c608] LATENCY=0
     -- Inputs
     layer0_node51_MUX_bit_math_h_l579_c3_c608_cond <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_cond;
     layer0_node51_MUX_bit_math_h_l579_c3_c608_iftrue <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_iftrue;
     layer0_node51_MUX_bit_math_h_l579_c3_c608_iffalse <= VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_iffalse;
     -- Outputs
     VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_return_output := layer0_node51_MUX_bit_math_h_l579_c3_c608_return_output;

     -- layer0_node8_MUX[bit_math_h_l106_c3_22f1] LATENCY=0
     -- Inputs
     layer0_node8_MUX_bit_math_h_l106_c3_22f1_cond <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_cond;
     layer0_node8_MUX_bit_math_h_l106_c3_22f1_iftrue <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_iftrue;
     layer0_node8_MUX_bit_math_h_l106_c3_22f1_iffalse <= VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_iffalse;
     -- Outputs
     VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_return_output := layer0_node8_MUX_bit_math_h_l106_c3_22f1_return_output;

     -- layer0_node20_MUX[bit_math_h_l238_c3_a0ec] LATENCY=0
     -- Inputs
     layer0_node20_MUX_bit_math_h_l238_c3_a0ec_cond <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_cond;
     layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iftrue <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iftrue;
     layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iffalse <= VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_iffalse;
     -- Outputs
     VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_return_output := layer0_node20_MUX_bit_math_h_l238_c3_a0ec_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_c2e4] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_c2e4_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_return_output := layer0_node7_MUX_bit_math_h_l95_c3_c2e4_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_2eec] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_2eec_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_2eec_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_2eec_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_return_output := layer0_node4_MUX_bit_math_h_l62_c3_2eec_return_output;

     -- layer0_node14_MUX[bit_math_h_l172_c3_e31d] LATENCY=0
     -- Inputs
     layer0_node14_MUX_bit_math_h_l172_c3_e31d_cond <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_cond;
     layer0_node14_MUX_bit_math_h_l172_c3_e31d_iftrue <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_iftrue;
     layer0_node14_MUX_bit_math_h_l172_c3_e31d_iffalse <= VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_iffalse;
     -- Outputs
     VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_return_output := layer0_node14_MUX_bit_math_h_l172_c3_e31d_return_output;

     -- layer0_node45_MUX[bit_math_h_l513_c3_1806] LATENCY=0
     -- Inputs
     layer0_node45_MUX_bit_math_h_l513_c3_1806_cond <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_cond;
     layer0_node45_MUX_bit_math_h_l513_c3_1806_iftrue <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_iftrue;
     layer0_node45_MUX_bit_math_h_l513_c3_1806_iffalse <= VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_iffalse;
     -- Outputs
     VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_return_output := layer0_node45_MUX_bit_math_h_l513_c3_1806_return_output;

     -- layer0_node35_MUX[bit_math_h_l403_c3_37e5] LATENCY=0
     -- Inputs
     layer0_node35_MUX_bit_math_h_l403_c3_37e5_cond <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_cond;
     layer0_node35_MUX_bit_math_h_l403_c3_37e5_iftrue <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_iftrue;
     layer0_node35_MUX_bit_math_h_l403_c3_37e5_iffalse <= VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_iffalse;
     -- Outputs
     VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_return_output := layer0_node35_MUX_bit_math_h_l403_c3_37e5_return_output;

     -- layer0_node6_MUX[bit_math_h_l84_c3_62aa] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_62aa_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_62aa_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_62aa_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_return_output := layer0_node6_MUX_bit_math_h_l84_c3_62aa_return_output;

     -- layer0_node23_MUX[bit_math_h_l271_c3_b2cd] LATENCY=0
     -- Inputs
     layer0_node23_MUX_bit_math_h_l271_c3_b2cd_cond <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_cond;
     layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iftrue <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iftrue;
     layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iffalse <= VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_iffalse;
     -- Outputs
     VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_return_output := layer0_node23_MUX_bit_math_h_l271_c3_b2cd_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_a274] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_a274_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_a274_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_a274_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_return_output := layer0_node3_MUX_bit_math_h_l51_c3_a274_return_output;

     -- layer0_node38_MUX[bit_math_h_l436_c3_b87e] LATENCY=0
     -- Inputs
     layer0_node38_MUX_bit_math_h_l436_c3_b87e_cond <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_cond;
     layer0_node38_MUX_bit_math_h_l436_c3_b87e_iftrue <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_iftrue;
     layer0_node38_MUX_bit_math_h_l436_c3_b87e_iffalse <= VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_iffalse;
     -- Outputs
     VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_return_output := layer0_node38_MUX_bit_math_h_l436_c3_b87e_return_output;

     -- layer0_node50_MUX[bit_math_h_l568_c3_ac6c] LATENCY=0
     -- Inputs
     layer0_node50_MUX_bit_math_h_l568_c3_ac6c_cond <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_cond;
     layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iftrue <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iftrue;
     layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iffalse <= VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_iffalse;
     -- Outputs
     VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_return_output := layer0_node50_MUX_bit_math_h_l568_c3_ac6c_return_output;

     -- layer0_node56_MUX[bit_math_h_l634_c3_259e] LATENCY=0
     -- Inputs
     layer0_node56_MUX_bit_math_h_l634_c3_259e_cond <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_cond;
     layer0_node56_MUX_bit_math_h_l634_c3_259e_iftrue <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_iftrue;
     layer0_node56_MUX_bit_math_h_l634_c3_259e_iffalse <= VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_iffalse;
     -- Outputs
     VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_return_output := layer0_node56_MUX_bit_math_h_l634_c3_259e_return_output;

     -- layer0_node27_MUX[bit_math_h_l315_c3_a6a8] LATENCY=0
     -- Inputs
     layer0_node27_MUX_bit_math_h_l315_c3_a6a8_cond <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_cond;
     layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iftrue <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iftrue;
     layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iffalse <= VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_iffalse;
     -- Outputs
     VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_return_output := layer0_node27_MUX_bit_math_h_l315_c3_a6a8_return_output;

     -- layer0_node54_MUX[bit_math_h_l612_c3_21f7] LATENCY=0
     -- Inputs
     layer0_node54_MUX_bit_math_h_l612_c3_21f7_cond <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_cond;
     layer0_node54_MUX_bit_math_h_l612_c3_21f7_iftrue <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_iftrue;
     layer0_node54_MUX_bit_math_h_l612_c3_21f7_iffalse <= VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_iffalse;
     -- Outputs
     VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_return_output := layer0_node54_MUX_bit_math_h_l612_c3_21f7_return_output;

     -- layer0_node32_MUX[bit_math_h_l370_c3_45be] LATENCY=0
     -- Inputs
     layer0_node32_MUX_bit_math_h_l370_c3_45be_cond <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_cond;
     layer0_node32_MUX_bit_math_h_l370_c3_45be_iftrue <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_iftrue;
     layer0_node32_MUX_bit_math_h_l370_c3_45be_iffalse <= VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_iffalse;
     -- Outputs
     VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_return_output := layer0_node32_MUX_bit_math_h_l370_c3_45be_return_output;

     -- layer0_node34_MUX[bit_math_h_l392_c3_7b48] LATENCY=0
     -- Inputs
     layer0_node34_MUX_bit_math_h_l392_c3_7b48_cond <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_cond;
     layer0_node34_MUX_bit_math_h_l392_c3_7b48_iftrue <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_iftrue;
     layer0_node34_MUX_bit_math_h_l392_c3_7b48_iffalse <= VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_iffalse;
     -- Outputs
     VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_return_output := layer0_node34_MUX_bit_math_h_l392_c3_7b48_return_output;

     -- layer0_node17_MUX[bit_math_h_l205_c3_ec06] LATENCY=0
     -- Inputs
     layer0_node17_MUX_bit_math_h_l205_c3_ec06_cond <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_cond;
     layer0_node17_MUX_bit_math_h_l205_c3_ec06_iftrue <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_iftrue;
     layer0_node17_MUX_bit_math_h_l205_c3_ec06_iffalse <= VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_iffalse;
     -- Outputs
     VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_return_output := layer0_node17_MUX_bit_math_h_l205_c3_ec06_return_output;

     -- layer0_node46_MUX[bit_math_h_l524_c3_c07c] LATENCY=0
     -- Inputs
     layer0_node46_MUX_bit_math_h_l524_c3_c07c_cond <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_cond;
     layer0_node46_MUX_bit_math_h_l524_c3_c07c_iftrue <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_iftrue;
     layer0_node46_MUX_bit_math_h_l524_c3_c07c_iffalse <= VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_iffalse;
     -- Outputs
     VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_return_output := layer0_node46_MUX_bit_math_h_l524_c3_c07c_return_output;

     -- layer0_node47_MUX[bit_math_h_l535_c3_a2fb] LATENCY=0
     -- Inputs
     layer0_node47_MUX_bit_math_h_l535_c3_a2fb_cond <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_cond;
     layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iftrue <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iftrue;
     layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iffalse <= VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_iffalse;
     -- Outputs
     VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_return_output := layer0_node47_MUX_bit_math_h_l535_c3_a2fb_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_85c1] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_85c1_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_85c1_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_85c1_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_return_output := layer0_node0_MUX_bit_math_h_l18_c3_85c1_return_output;

     -- layer0_node29_MUX[bit_math_h_l337_c3_1d84] LATENCY=0
     -- Inputs
     layer0_node29_MUX_bit_math_h_l337_c3_1d84_cond <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_cond;
     layer0_node29_MUX_bit_math_h_l337_c3_1d84_iftrue <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_iftrue;
     layer0_node29_MUX_bit_math_h_l337_c3_1d84_iffalse <= VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_iffalse;
     -- Outputs
     VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_return_output := layer0_node29_MUX_bit_math_h_l337_c3_1d84_return_output;

     -- layer0_node19_MUX[bit_math_h_l227_c3_0da7] LATENCY=0
     -- Inputs
     layer0_node19_MUX_bit_math_h_l227_c3_0da7_cond <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_cond;
     layer0_node19_MUX_bit_math_h_l227_c3_0da7_iftrue <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_iftrue;
     layer0_node19_MUX_bit_math_h_l227_c3_0da7_iffalse <= VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_iffalse;
     -- Outputs
     VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_return_output := layer0_node19_MUX_bit_math_h_l227_c3_0da7_return_output;

     -- layer0_node59_MUX[bit_math_h_l667_c3_060a] LATENCY=0
     -- Inputs
     layer0_node59_MUX_bit_math_h_l667_c3_060a_cond <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_cond;
     layer0_node59_MUX_bit_math_h_l667_c3_060a_iftrue <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_iftrue;
     layer0_node59_MUX_bit_math_h_l667_c3_060a_iffalse <= VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_iffalse;
     -- Outputs
     VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_return_output := layer0_node59_MUX_bit_math_h_l667_c3_060a_return_output;

     -- layer0_node18_MUX[bit_math_h_l216_c3_7962] LATENCY=0
     -- Inputs
     layer0_node18_MUX_bit_math_h_l216_c3_7962_cond <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_cond;
     layer0_node18_MUX_bit_math_h_l216_c3_7962_iftrue <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_iftrue;
     layer0_node18_MUX_bit_math_h_l216_c3_7962_iffalse <= VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_iffalse;
     -- Outputs
     VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_return_output := layer0_node18_MUX_bit_math_h_l216_c3_7962_return_output;

     -- layer0_node9_MUX[bit_math_h_l117_c3_391b] LATENCY=0
     -- Inputs
     layer0_node9_MUX_bit_math_h_l117_c3_391b_cond <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_cond;
     layer0_node9_MUX_bit_math_h_l117_c3_391b_iftrue <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_iftrue;
     layer0_node9_MUX_bit_math_h_l117_c3_391b_iffalse <= VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_iffalse;
     -- Outputs
     VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_return_output := layer0_node9_MUX_bit_math_h_l117_c3_391b_return_output;

     -- layer0_node55_MUX[bit_math_h_l623_c3_a654] LATENCY=0
     -- Inputs
     layer0_node55_MUX_bit_math_h_l623_c3_a654_cond <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_cond;
     layer0_node55_MUX_bit_math_h_l623_c3_a654_iftrue <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_iftrue;
     layer0_node55_MUX_bit_math_h_l623_c3_a654_iffalse <= VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_iffalse;
     -- Outputs
     VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_return_output := layer0_node55_MUX_bit_math_h_l623_c3_a654_return_output;

     -- layer0_node5_MUX[bit_math_h_l73_c3_5736] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_5736_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_5736_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_5736_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_return_output := layer0_node5_MUX_bit_math_h_l73_c3_5736_return_output;

     -- layer0_node52_MUX[bit_math_h_l590_c3_f975] LATENCY=0
     -- Inputs
     layer0_node52_MUX_bit_math_h_l590_c3_f975_cond <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_cond;
     layer0_node52_MUX_bit_math_h_l590_c3_f975_iftrue <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_iftrue;
     layer0_node52_MUX_bit_math_h_l590_c3_f975_iffalse <= VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_iffalse;
     -- Outputs
     VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_return_output := layer0_node52_MUX_bit_math_h_l590_c3_f975_return_output;

     -- layer0_node15_MUX[bit_math_h_l183_c3_313e] LATENCY=0
     -- Inputs
     layer0_node15_MUX_bit_math_h_l183_c3_313e_cond <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_cond;
     layer0_node15_MUX_bit_math_h_l183_c3_313e_iftrue <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_iftrue;
     layer0_node15_MUX_bit_math_h_l183_c3_313e_iffalse <= VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_iffalse;
     -- Outputs
     VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_return_output := layer0_node15_MUX_bit_math_h_l183_c3_313e_return_output;

     -- layer0_node60_MUX[bit_math_h_l678_c3_dedf] LATENCY=0
     -- Inputs
     layer0_node60_MUX_bit_math_h_l678_c3_dedf_cond <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_cond;
     layer0_node60_MUX_bit_math_h_l678_c3_dedf_iftrue <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_iftrue;
     layer0_node60_MUX_bit_math_h_l678_c3_dedf_iffalse <= VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_iffalse;
     -- Outputs
     VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_return_output := layer0_node60_MUX_bit_math_h_l678_c3_dedf_return_output;

     -- layer0_node33_MUX[bit_math_h_l381_c3_2a50] LATENCY=0
     -- Inputs
     layer0_node33_MUX_bit_math_h_l381_c3_2a50_cond <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_cond;
     layer0_node33_MUX_bit_math_h_l381_c3_2a50_iftrue <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_iftrue;
     layer0_node33_MUX_bit_math_h_l381_c3_2a50_iffalse <= VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_iffalse;
     -- Outputs
     VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_return_output := layer0_node33_MUX_bit_math_h_l381_c3_2a50_return_output;

     -- layer0_node43_MUX[bit_math_h_l491_c3_a5e9] LATENCY=0
     -- Inputs
     layer0_node43_MUX_bit_math_h_l491_c3_a5e9_cond <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_cond;
     layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iftrue <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iftrue;
     layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iffalse <= VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_iffalse;
     -- Outputs
     VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_return_output := layer0_node43_MUX_bit_math_h_l491_c3_a5e9_return_output;

     -- layer0_node40_MUX[bit_math_h_l458_c3_a82d] LATENCY=0
     -- Inputs
     layer0_node40_MUX_bit_math_h_l458_c3_a82d_cond <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_cond;
     layer0_node40_MUX_bit_math_h_l458_c3_a82d_iftrue <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_iftrue;
     layer0_node40_MUX_bit_math_h_l458_c3_a82d_iffalse <= VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_iffalse;
     -- Outputs
     VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_return_output := layer0_node40_MUX_bit_math_h_l458_c3_a82d_return_output;

     -- layer0_node22_MUX[bit_math_h_l260_c3_50aa] LATENCY=0
     -- Inputs
     layer0_node22_MUX_bit_math_h_l260_c3_50aa_cond <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_cond;
     layer0_node22_MUX_bit_math_h_l260_c3_50aa_iftrue <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_iftrue;
     layer0_node22_MUX_bit_math_h_l260_c3_50aa_iffalse <= VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_iffalse;
     -- Outputs
     VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_return_output := layer0_node22_MUX_bit_math_h_l260_c3_50aa_return_output;

     -- layer0_node49_MUX[bit_math_h_l557_c3_5e53] LATENCY=0
     -- Inputs
     layer0_node49_MUX_bit_math_h_l557_c3_5e53_cond <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_cond;
     layer0_node49_MUX_bit_math_h_l557_c3_5e53_iftrue <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_iftrue;
     layer0_node49_MUX_bit_math_h_l557_c3_5e53_iffalse <= VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_iffalse;
     -- Outputs
     VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_return_output := layer0_node49_MUX_bit_math_h_l557_c3_5e53_return_output;

     -- layer0_node62_MUX[bit_math_h_l700_c3_7046] LATENCY=0
     -- Inputs
     layer0_node62_MUX_bit_math_h_l700_c3_7046_cond <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_cond;
     layer0_node62_MUX_bit_math_h_l700_c3_7046_iftrue <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_iftrue;
     layer0_node62_MUX_bit_math_h_l700_c3_7046_iffalse <= VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_iffalse;
     -- Outputs
     VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_return_output := layer0_node62_MUX_bit_math_h_l700_c3_7046_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_43b7] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_43b7_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_43b7_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_43b7_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_return_output := layer0_node2_MUX_bit_math_h_l40_c3_43b7_return_output;

     -- layer0_node26_MUX[bit_math_h_l304_c3_809a] LATENCY=0
     -- Inputs
     layer0_node26_MUX_bit_math_h_l304_c3_809a_cond <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_cond;
     layer0_node26_MUX_bit_math_h_l304_c3_809a_iftrue <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_iftrue;
     layer0_node26_MUX_bit_math_h_l304_c3_809a_iffalse <= VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_iffalse;
     -- Outputs
     VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_return_output := layer0_node26_MUX_bit_math_h_l304_c3_809a_return_output;

     -- layer0_node25_MUX[bit_math_h_l293_c3_d8bb] LATENCY=0
     -- Inputs
     layer0_node25_MUX_bit_math_h_l293_c3_d8bb_cond <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_cond;
     layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iftrue <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iftrue;
     layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iffalse <= VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_iffalse;
     -- Outputs
     VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_return_output := layer0_node25_MUX_bit_math_h_l293_c3_d8bb_return_output;

     -- layer0_node24_MUX[bit_math_h_l282_c3_0847] LATENCY=0
     -- Inputs
     layer0_node24_MUX_bit_math_h_l282_c3_0847_cond <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_cond;
     layer0_node24_MUX_bit_math_h_l282_c3_0847_iftrue <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_iftrue;
     layer0_node24_MUX_bit_math_h_l282_c3_0847_iffalse <= VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_iffalse;
     -- Outputs
     VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_return_output := layer0_node24_MUX_bit_math_h_l282_c3_0847_return_output;

     -- layer0_node44_MUX[bit_math_h_l502_c3_7ff6] LATENCY=0
     -- Inputs
     layer0_node44_MUX_bit_math_h_l502_c3_7ff6_cond <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_cond;
     layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iftrue <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iftrue;
     layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iffalse <= VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_iffalse;
     -- Outputs
     VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_return_output := layer0_node44_MUX_bit_math_h_l502_c3_7ff6_return_output;

     -- layer0_node53_MUX[bit_math_h_l601_c3_86a8] LATENCY=0
     -- Inputs
     layer0_node53_MUX_bit_math_h_l601_c3_86a8_cond <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_cond;
     layer0_node53_MUX_bit_math_h_l601_c3_86a8_iftrue <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_iftrue;
     layer0_node53_MUX_bit_math_h_l601_c3_86a8_iffalse <= VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_iffalse;
     -- Outputs
     VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_return_output := layer0_node53_MUX_bit_math_h_l601_c3_86a8_return_output;

     -- layer0_node30_MUX[bit_math_h_l348_c3_27f8] LATENCY=0
     -- Inputs
     layer0_node30_MUX_bit_math_h_l348_c3_27f8_cond <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_cond;
     layer0_node30_MUX_bit_math_h_l348_c3_27f8_iftrue <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_iftrue;
     layer0_node30_MUX_bit_math_h_l348_c3_27f8_iffalse <= VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_iffalse;
     -- Outputs
     VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_return_output := layer0_node30_MUX_bit_math_h_l348_c3_27f8_return_output;

     -- layer0_node31_MUX[bit_math_h_l359_c3_e962] LATENCY=0
     -- Inputs
     layer0_node31_MUX_bit_math_h_l359_c3_e962_cond <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_cond;
     layer0_node31_MUX_bit_math_h_l359_c3_e962_iftrue <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_iftrue;
     layer0_node31_MUX_bit_math_h_l359_c3_e962_iffalse <= VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_iffalse;
     -- Outputs
     VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_return_output := layer0_node31_MUX_bit_math_h_l359_c3_e962_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_85c1_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_iffalse := VAR_layer0_node10_MUX_bit_math_h_l128_c3_1e58_return_output;
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_iftrue := VAR_layer0_node11_MUX_bit_math_h_l139_c3_6d2d_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iffalse := VAR_layer0_node12_MUX_bit_math_h_l150_c3_40e1_return_output;
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iftrue := VAR_layer0_node13_MUX_bit_math_h_l161_c3_28f7_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_iffalse := VAR_layer0_node14_MUX_bit_math_h_l172_c3_e31d_return_output;
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_iftrue := VAR_layer0_node15_MUX_bit_math_h_l183_c3_313e_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_iffalse := VAR_layer0_node16_MUX_bit_math_h_l194_c3_614a_return_output;
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_iftrue := VAR_layer0_node17_MUX_bit_math_h_l205_c3_ec06_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_iffalse := VAR_layer0_node18_MUX_bit_math_h_l216_c3_7962_return_output;
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_iftrue := VAR_layer0_node19_MUX_bit_math_h_l227_c3_0da7_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_a7d4_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iffalse := VAR_layer0_node20_MUX_bit_math_h_l238_c3_a0ec_return_output;
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iftrue := VAR_layer0_node21_MUX_bit_math_h_l249_c3_a3f0_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_iffalse := VAR_layer0_node22_MUX_bit_math_h_l260_c3_50aa_return_output;
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_iftrue := VAR_layer0_node23_MUX_bit_math_h_l271_c3_b2cd_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_iffalse := VAR_layer0_node24_MUX_bit_math_h_l282_c3_0847_return_output;
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_iftrue := VAR_layer0_node25_MUX_bit_math_h_l293_c3_d8bb_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iffalse := VAR_layer0_node26_MUX_bit_math_h_l304_c3_809a_return_output;
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iftrue := VAR_layer0_node27_MUX_bit_math_h_l315_c3_a6a8_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_iffalse := VAR_layer0_node28_MUX_bit_math_h_l326_c3_b62d_return_output;
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_iftrue := VAR_layer0_node29_MUX_bit_math_h_l337_c3_1d84_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_43b7_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_iffalse := VAR_layer0_node30_MUX_bit_math_h_l348_c3_27f8_return_output;
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_iftrue := VAR_layer0_node31_MUX_bit_math_h_l359_c3_e962_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iffalse := VAR_layer0_node32_MUX_bit_math_h_l370_c3_45be_return_output;
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iftrue := VAR_layer0_node33_MUX_bit_math_h_l381_c3_2a50_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iffalse := VAR_layer0_node34_MUX_bit_math_h_l392_c3_7b48_return_output;
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iftrue := VAR_layer0_node35_MUX_bit_math_h_l403_c3_37e5_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_iffalse := VAR_layer0_node36_MUX_bit_math_h_l414_c3_fd1a_return_output;
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_iftrue := VAR_layer0_node37_MUX_bit_math_h_l425_c3_8edb_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_iffalse := VAR_layer0_node38_MUX_bit_math_h_l436_c3_b87e_return_output;
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_iftrue := VAR_layer0_node39_MUX_bit_math_h_l447_c3_8780_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_a274_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_iffalse := VAR_layer0_node40_MUX_bit_math_h_l458_c3_a82d_return_output;
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_iftrue := VAR_layer0_node41_MUX_bit_math_h_l469_c3_f332_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_iffalse := VAR_layer0_node42_MUX_bit_math_h_l480_c3_8296_return_output;
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_iftrue := VAR_layer0_node43_MUX_bit_math_h_l491_c3_a5e9_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_iffalse := VAR_layer0_node44_MUX_bit_math_h_l502_c3_7ff6_return_output;
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_iftrue := VAR_layer0_node45_MUX_bit_math_h_l513_c3_1806_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_iffalse := VAR_layer0_node46_MUX_bit_math_h_l524_c3_c07c_return_output;
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_iftrue := VAR_layer0_node47_MUX_bit_math_h_l535_c3_a2fb_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iffalse := VAR_layer0_node48_MUX_bit_math_h_l546_c3_a700_return_output;
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iftrue := VAR_layer0_node49_MUX_bit_math_h_l557_c3_5e53_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_2eec_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iffalse := VAR_layer0_node50_MUX_bit_math_h_l568_c3_ac6c_return_output;
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iftrue := VAR_layer0_node51_MUX_bit_math_h_l579_c3_c608_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iffalse := VAR_layer0_node52_MUX_bit_math_h_l590_c3_f975_return_output;
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iftrue := VAR_layer0_node53_MUX_bit_math_h_l601_c3_86a8_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_iffalse := VAR_layer0_node54_MUX_bit_math_h_l612_c3_21f7_return_output;
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_iftrue := VAR_layer0_node55_MUX_bit_math_h_l623_c3_a654_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_iffalse := VAR_layer0_node56_MUX_bit_math_h_l634_c3_259e_return_output;
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_iftrue := VAR_layer0_node57_MUX_bit_math_h_l645_c3_3acf_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iffalse := VAR_layer0_node58_MUX_bit_math_h_l656_c3_6a0d_return_output;
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iftrue := VAR_layer0_node59_MUX_bit_math_h_l667_c3_060a_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_5736_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iffalse := VAR_layer0_node60_MUX_bit_math_h_l678_c3_dedf_return_output;
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iftrue := VAR_layer0_node61_MUX_bit_math_h_l689_c3_26a3_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_iffalse := VAR_layer0_node62_MUX_bit_math_h_l700_c3_7046_return_output;
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_iftrue := VAR_layer0_node63_MUX_bit_math_h_l711_c3_0125_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_62aa_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_c2e4_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_iffalse := VAR_layer0_node8_MUX_bit_math_h_l106_c3_22f1_return_output;
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_iftrue := VAR_layer0_node9_MUX_bit_math_h_l117_c3_391b_return_output;
     -- layer1_node12_MUX[bit_math_h_l860_c3_7af8] LATENCY=0
     -- Inputs
     layer1_node12_MUX_bit_math_h_l860_c3_7af8_cond <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_cond;
     layer1_node12_MUX_bit_math_h_l860_c3_7af8_iftrue <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_iftrue;
     layer1_node12_MUX_bit_math_h_l860_c3_7af8_iffalse <= VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_iffalse;
     -- Outputs
     VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_return_output := layer1_node12_MUX_bit_math_h_l860_c3_7af8_return_output;

     -- layer1_node28_MUX[bit_math_h_l1036_c3_f568] LATENCY=0
     -- Inputs
     layer1_node28_MUX_bit_math_h_l1036_c3_f568_cond <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_cond;
     layer1_node28_MUX_bit_math_h_l1036_c3_f568_iftrue <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_iftrue;
     layer1_node28_MUX_bit_math_h_l1036_c3_f568_iffalse <= VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_iffalse;
     -- Outputs
     VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_return_output := layer1_node28_MUX_bit_math_h_l1036_c3_f568_return_output;

     -- layer1_node3_MUX[bit_math_h_l761_c3_123f] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l761_c3_123f_cond <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_cond;
     layer1_node3_MUX_bit_math_h_l761_c3_123f_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_iftrue;
     layer1_node3_MUX_bit_math_h_l761_c3_123f_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_return_output := layer1_node3_MUX_bit_math_h_l761_c3_123f_return_output;

     -- layer1_node15_MUX[bit_math_h_l893_c3_3f51] LATENCY=0
     -- Inputs
     layer1_node15_MUX_bit_math_h_l893_c3_3f51_cond <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_cond;
     layer1_node15_MUX_bit_math_h_l893_c3_3f51_iftrue <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_iftrue;
     layer1_node15_MUX_bit_math_h_l893_c3_3f51_iffalse <= VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_iffalse;
     -- Outputs
     VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_return_output := layer1_node15_MUX_bit_math_h_l893_c3_3f51_return_output;

     -- layer1_node18_MUX[bit_math_h_l926_c3_5844] LATENCY=0
     -- Inputs
     layer1_node18_MUX_bit_math_h_l926_c3_5844_cond <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_cond;
     layer1_node18_MUX_bit_math_h_l926_c3_5844_iftrue <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_iftrue;
     layer1_node18_MUX_bit_math_h_l926_c3_5844_iffalse <= VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_iffalse;
     -- Outputs
     VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_return_output := layer1_node18_MUX_bit_math_h_l926_c3_5844_return_output;

     -- layer1_node19_MUX[bit_math_h_l937_c3_7dba] LATENCY=0
     -- Inputs
     layer1_node19_MUX_bit_math_h_l937_c3_7dba_cond <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_cond;
     layer1_node19_MUX_bit_math_h_l937_c3_7dba_iftrue <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_iftrue;
     layer1_node19_MUX_bit_math_h_l937_c3_7dba_iffalse <= VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_iffalse;
     -- Outputs
     VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_return_output := layer1_node19_MUX_bit_math_h_l937_c3_7dba_return_output;

     -- layer1_node22_MUX[bit_math_h_l970_c3_65bd] LATENCY=0
     -- Inputs
     layer1_node22_MUX_bit_math_h_l970_c3_65bd_cond <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_cond;
     layer1_node22_MUX_bit_math_h_l970_c3_65bd_iftrue <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_iftrue;
     layer1_node22_MUX_bit_math_h_l970_c3_65bd_iffalse <= VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_iffalse;
     -- Outputs
     VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_return_output := layer1_node22_MUX_bit_math_h_l970_c3_65bd_return_output;

     -- layer1_node31_MUX[bit_math_h_l1069_c3_6881] LATENCY=0
     -- Inputs
     layer1_node31_MUX_bit_math_h_l1069_c3_6881_cond <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_cond;
     layer1_node31_MUX_bit_math_h_l1069_c3_6881_iftrue <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_iftrue;
     layer1_node31_MUX_bit_math_h_l1069_c3_6881_iffalse <= VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_iffalse;
     -- Outputs
     VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_return_output := layer1_node31_MUX_bit_math_h_l1069_c3_6881_return_output;

     -- layer1_node24_MUX[bit_math_h_l992_c3_8ee7] LATENCY=0
     -- Inputs
     layer1_node24_MUX_bit_math_h_l992_c3_8ee7_cond <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_cond;
     layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iftrue <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iftrue;
     layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iffalse <= VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_iffalse;
     -- Outputs
     VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_return_output := layer1_node24_MUX_bit_math_h_l992_c3_8ee7_return_output;

     -- layer1_node5_MUX[bit_math_h_l783_c3_58a8] LATENCY=0
     -- Inputs
     layer1_node5_MUX_bit_math_h_l783_c3_58a8_cond <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_cond;
     layer1_node5_MUX_bit_math_h_l783_c3_58a8_iftrue <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_iftrue;
     layer1_node5_MUX_bit_math_h_l783_c3_58a8_iffalse <= VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_iffalse;
     -- Outputs
     VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_return_output := layer1_node5_MUX_bit_math_h_l783_c3_58a8_return_output;

     -- layer1_node2_MUX[bit_math_h_l750_c3_e4a0] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l750_c3_e4a0_cond <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_cond;
     layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iftrue;
     layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_return_output := layer1_node2_MUX_bit_math_h_l750_c3_e4a0_return_output;

     -- layer1_node16_MUX[bit_math_h_l904_c3_e9a5] LATENCY=0
     -- Inputs
     layer1_node16_MUX_bit_math_h_l904_c3_e9a5_cond <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_cond;
     layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iftrue <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iftrue;
     layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iffalse <= VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_iffalse;
     -- Outputs
     VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_return_output := layer1_node16_MUX_bit_math_h_l904_c3_e9a5_return_output;

     -- layer1_node27_MUX[bit_math_h_l1025_c3_465f] LATENCY=0
     -- Inputs
     layer1_node27_MUX_bit_math_h_l1025_c3_465f_cond <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_cond;
     layer1_node27_MUX_bit_math_h_l1025_c3_465f_iftrue <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_iftrue;
     layer1_node27_MUX_bit_math_h_l1025_c3_465f_iffalse <= VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_iffalse;
     -- Outputs
     VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_return_output := layer1_node27_MUX_bit_math_h_l1025_c3_465f_return_output;

     -- layer1_node0_MUX[bit_math_h_l728_c3_287e] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l728_c3_287e_cond <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_cond;
     layer1_node0_MUX_bit_math_h_l728_c3_287e_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_iftrue;
     layer1_node0_MUX_bit_math_h_l728_c3_287e_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_return_output := layer1_node0_MUX_bit_math_h_l728_c3_287e_return_output;

     -- layer1_node1_MUX[bit_math_h_l739_c3_3eb3] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l739_c3_3eb3_cond <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_cond;
     layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iftrue;
     layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_return_output := layer1_node1_MUX_bit_math_h_l739_c3_3eb3_return_output;

     -- layer1_node14_MUX[bit_math_h_l882_c3_10cf] LATENCY=0
     -- Inputs
     layer1_node14_MUX_bit_math_h_l882_c3_10cf_cond <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_cond;
     layer1_node14_MUX_bit_math_h_l882_c3_10cf_iftrue <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_iftrue;
     layer1_node14_MUX_bit_math_h_l882_c3_10cf_iffalse <= VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_iffalse;
     -- Outputs
     VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_return_output := layer1_node14_MUX_bit_math_h_l882_c3_10cf_return_output;

     -- layer1_node26_MUX[bit_math_h_l1014_c3_d8aa] LATENCY=0
     -- Inputs
     layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_cond <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_cond;
     layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iftrue <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iftrue;
     layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iffalse <= VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_iffalse;
     -- Outputs
     VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_return_output := layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_return_output;

     -- layer1_node20_MUX[bit_math_h_l948_c3_2725] LATENCY=0
     -- Inputs
     layer1_node20_MUX_bit_math_h_l948_c3_2725_cond <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_cond;
     layer1_node20_MUX_bit_math_h_l948_c3_2725_iftrue <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_iftrue;
     layer1_node20_MUX_bit_math_h_l948_c3_2725_iffalse <= VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_iffalse;
     -- Outputs
     VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_return_output := layer1_node20_MUX_bit_math_h_l948_c3_2725_return_output;

     -- layer1_node8_MUX[bit_math_h_l816_c3_db42] LATENCY=0
     -- Inputs
     layer1_node8_MUX_bit_math_h_l816_c3_db42_cond <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_cond;
     layer1_node8_MUX_bit_math_h_l816_c3_db42_iftrue <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_iftrue;
     layer1_node8_MUX_bit_math_h_l816_c3_db42_iffalse <= VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_iffalse;
     -- Outputs
     VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_return_output := layer1_node8_MUX_bit_math_h_l816_c3_db42_return_output;

     -- layer1_node29_MUX[bit_math_h_l1047_c3_8f77] LATENCY=0
     -- Inputs
     layer1_node29_MUX_bit_math_h_l1047_c3_8f77_cond <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_cond;
     layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iftrue <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iftrue;
     layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iffalse <= VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_iffalse;
     -- Outputs
     VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_return_output := layer1_node29_MUX_bit_math_h_l1047_c3_8f77_return_output;

     -- layer1_node10_MUX[bit_math_h_l838_c3_a2e2] LATENCY=0
     -- Inputs
     layer1_node10_MUX_bit_math_h_l838_c3_a2e2_cond <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_cond;
     layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iftrue <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iftrue;
     layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iffalse <= VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_iffalse;
     -- Outputs
     VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_return_output := layer1_node10_MUX_bit_math_h_l838_c3_a2e2_return_output;

     -- layer1_node4_MUX[bit_math_h_l772_c3_0289] LATENCY=0
     -- Inputs
     layer1_node4_MUX_bit_math_h_l772_c3_0289_cond <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_cond;
     layer1_node4_MUX_bit_math_h_l772_c3_0289_iftrue <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_iftrue;
     layer1_node4_MUX_bit_math_h_l772_c3_0289_iffalse <= VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_iffalse;
     -- Outputs
     VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_return_output := layer1_node4_MUX_bit_math_h_l772_c3_0289_return_output;

     -- layer1_node21_MUX[bit_math_h_l959_c3_8499] LATENCY=0
     -- Inputs
     layer1_node21_MUX_bit_math_h_l959_c3_8499_cond <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_cond;
     layer1_node21_MUX_bit_math_h_l959_c3_8499_iftrue <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_iftrue;
     layer1_node21_MUX_bit_math_h_l959_c3_8499_iffalse <= VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_iffalse;
     -- Outputs
     VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_return_output := layer1_node21_MUX_bit_math_h_l959_c3_8499_return_output;

     -- layer1_node7_MUX[bit_math_h_l805_c3_1224] LATENCY=0
     -- Inputs
     layer1_node7_MUX_bit_math_h_l805_c3_1224_cond <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_cond;
     layer1_node7_MUX_bit_math_h_l805_c3_1224_iftrue <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_iftrue;
     layer1_node7_MUX_bit_math_h_l805_c3_1224_iffalse <= VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_iffalse;
     -- Outputs
     VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_return_output := layer1_node7_MUX_bit_math_h_l805_c3_1224_return_output;

     -- layer1_node6_MUX[bit_math_h_l794_c3_ebf4] LATENCY=0
     -- Inputs
     layer1_node6_MUX_bit_math_h_l794_c3_ebf4_cond <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_cond;
     layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iftrue <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iftrue;
     layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iffalse <= VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_iffalse;
     -- Outputs
     VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_return_output := layer1_node6_MUX_bit_math_h_l794_c3_ebf4_return_output;

     -- layer1_node23_MUX[bit_math_h_l981_c3_3335] LATENCY=0
     -- Inputs
     layer1_node23_MUX_bit_math_h_l981_c3_3335_cond <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_cond;
     layer1_node23_MUX_bit_math_h_l981_c3_3335_iftrue <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_iftrue;
     layer1_node23_MUX_bit_math_h_l981_c3_3335_iffalse <= VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_iffalse;
     -- Outputs
     VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_return_output := layer1_node23_MUX_bit_math_h_l981_c3_3335_return_output;

     -- layer1_node30_MUX[bit_math_h_l1058_c3_d4dc] LATENCY=0
     -- Inputs
     layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_cond <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_cond;
     layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iftrue <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iftrue;
     layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iffalse <= VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_iffalse;
     -- Outputs
     VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_return_output := layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_return_output;

     -- layer1_node9_MUX[bit_math_h_l827_c3_8290] LATENCY=0
     -- Inputs
     layer1_node9_MUX_bit_math_h_l827_c3_8290_cond <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_cond;
     layer1_node9_MUX_bit_math_h_l827_c3_8290_iftrue <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_iftrue;
     layer1_node9_MUX_bit_math_h_l827_c3_8290_iffalse <= VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_iffalse;
     -- Outputs
     VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_return_output := layer1_node9_MUX_bit_math_h_l827_c3_8290_return_output;

     -- layer1_node13_MUX[bit_math_h_l871_c3_d1fd] LATENCY=0
     -- Inputs
     layer1_node13_MUX_bit_math_h_l871_c3_d1fd_cond <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_cond;
     layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iftrue <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iftrue;
     layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iffalse <= VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_iffalse;
     -- Outputs
     VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_return_output := layer1_node13_MUX_bit_math_h_l871_c3_d1fd_return_output;

     -- layer1_node11_MUX[bit_math_h_l849_c3_dc54] LATENCY=0
     -- Inputs
     layer1_node11_MUX_bit_math_h_l849_c3_dc54_cond <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_cond;
     layer1_node11_MUX_bit_math_h_l849_c3_dc54_iftrue <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_iftrue;
     layer1_node11_MUX_bit_math_h_l849_c3_dc54_iffalse <= VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_iffalse;
     -- Outputs
     VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_return_output := layer1_node11_MUX_bit_math_h_l849_c3_dc54_return_output;

     -- layer1_node17_MUX[bit_math_h_l915_c3_4b4e] LATENCY=0
     -- Inputs
     layer1_node17_MUX_bit_math_h_l915_c3_4b4e_cond <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_cond;
     layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iftrue <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iftrue;
     layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iffalse <= VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_iffalse;
     -- Outputs
     VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_return_output := layer1_node17_MUX_bit_math_h_l915_c3_4b4e_return_output;

     -- layer1_node25_MUX[bit_math_h_l1003_c3_8e94] LATENCY=0
     -- Inputs
     layer1_node25_MUX_bit_math_h_l1003_c3_8e94_cond <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_cond;
     layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iftrue <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iftrue;
     layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iffalse <= VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_iffalse;
     -- Outputs
     VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_return_output := layer1_node25_MUX_bit_math_h_l1003_c3_8e94_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iffalse := VAR_layer1_node0_MUX_bit_math_h_l728_c3_287e_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_iffalse := VAR_layer1_node10_MUX_bit_math_h_l838_c3_a2e2_return_output;
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_iftrue := VAR_layer1_node11_MUX_bit_math_h_l849_c3_dc54_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_iffalse := VAR_layer1_node12_MUX_bit_math_h_l860_c3_7af8_return_output;
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_iftrue := VAR_layer1_node13_MUX_bit_math_h_l871_c3_d1fd_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_iffalse := VAR_layer1_node14_MUX_bit_math_h_l882_c3_10cf_return_output;
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_iftrue := VAR_layer1_node15_MUX_bit_math_h_l893_c3_3f51_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_iffalse := VAR_layer1_node16_MUX_bit_math_h_l904_c3_e9a5_return_output;
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_iftrue := VAR_layer1_node17_MUX_bit_math_h_l915_c3_4b4e_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iffalse := VAR_layer1_node18_MUX_bit_math_h_l926_c3_5844_return_output;
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iftrue := VAR_layer1_node19_MUX_bit_math_h_l937_c3_7dba_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iftrue := VAR_layer1_node1_MUX_bit_math_h_l739_c3_3eb3_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_iffalse := VAR_layer1_node20_MUX_bit_math_h_l948_c3_2725_return_output;
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_iftrue := VAR_layer1_node21_MUX_bit_math_h_l959_c3_8499_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iffalse := VAR_layer1_node22_MUX_bit_math_h_l970_c3_65bd_return_output;
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iftrue := VAR_layer1_node23_MUX_bit_math_h_l981_c3_3335_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iffalse := VAR_layer1_node24_MUX_bit_math_h_l992_c3_8ee7_return_output;
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iftrue := VAR_layer1_node25_MUX_bit_math_h_l1003_c3_8e94_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iffalse := VAR_layer1_node26_MUX_bit_math_h_l1014_c3_d8aa_return_output;
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iftrue := VAR_layer1_node27_MUX_bit_math_h_l1025_c3_465f_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iffalse := VAR_layer1_node28_MUX_bit_math_h_l1036_c3_f568_return_output;
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iftrue := VAR_layer1_node29_MUX_bit_math_h_l1047_c3_8f77_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iffalse := VAR_layer1_node2_MUX_bit_math_h_l750_c3_e4a0_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iffalse := VAR_layer1_node30_MUX_bit_math_h_l1058_c3_d4dc_return_output;
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iftrue := VAR_layer1_node31_MUX_bit_math_h_l1069_c3_6881_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iftrue := VAR_layer1_node3_MUX_bit_math_h_l761_c3_123f_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iffalse := VAR_layer1_node4_MUX_bit_math_h_l772_c3_0289_return_output;
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iftrue := VAR_layer1_node5_MUX_bit_math_h_l783_c3_58a8_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iffalse := VAR_layer1_node6_MUX_bit_math_h_l794_c3_ebf4_return_output;
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iftrue := VAR_layer1_node7_MUX_bit_math_h_l805_c3_1224_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iffalse := VAR_layer1_node8_MUX_bit_math_h_l816_c3_db42_return_output;
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iftrue := VAR_layer1_node9_MUX_bit_math_h_l827_c3_8290_return_output;
     -- layer2_node11_MUX[bit_math_h_l1207_c3_80d7] LATENCY=0
     -- Inputs
     layer2_node11_MUX_bit_math_h_l1207_c3_80d7_cond <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_cond;
     layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iftrue <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iftrue;
     layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iffalse <= VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_iffalse;
     -- Outputs
     VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_return_output := layer2_node11_MUX_bit_math_h_l1207_c3_80d7_return_output;

     -- layer2_node8_MUX[bit_math_h_l1174_c3_918c] LATENCY=0
     -- Inputs
     layer2_node8_MUX_bit_math_h_l1174_c3_918c_cond <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_cond;
     layer2_node8_MUX_bit_math_h_l1174_c3_918c_iftrue <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_iftrue;
     layer2_node8_MUX_bit_math_h_l1174_c3_918c_iffalse <= VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_iffalse;
     -- Outputs
     VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_return_output := layer2_node8_MUX_bit_math_h_l1174_c3_918c_return_output;

     -- layer2_node6_MUX[bit_math_h_l1152_c3_be62] LATENCY=0
     -- Inputs
     layer2_node6_MUX_bit_math_h_l1152_c3_be62_cond <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_cond;
     layer2_node6_MUX_bit_math_h_l1152_c3_be62_iftrue <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_iftrue;
     layer2_node6_MUX_bit_math_h_l1152_c3_be62_iffalse <= VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_iffalse;
     -- Outputs
     VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_return_output := layer2_node6_MUX_bit_math_h_l1152_c3_be62_return_output;

     -- layer2_node2_MUX[bit_math_h_l1108_c3_0b56] LATENCY=0
     -- Inputs
     layer2_node2_MUX_bit_math_h_l1108_c3_0b56_cond <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_cond;
     layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iftrue <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iftrue;
     layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iffalse <= VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_iffalse;
     -- Outputs
     VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_return_output := layer2_node2_MUX_bit_math_h_l1108_c3_0b56_return_output;

     -- layer2_node3_MUX[bit_math_h_l1119_c3_7df6] LATENCY=0
     -- Inputs
     layer2_node3_MUX_bit_math_h_l1119_c3_7df6_cond <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_cond;
     layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iftrue <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iftrue;
     layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iffalse <= VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_iffalse;
     -- Outputs
     VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_return_output := layer2_node3_MUX_bit_math_h_l1119_c3_7df6_return_output;

     -- layer2_node0_MUX[bit_math_h_l1086_c3_f1d8] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_cond <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_cond;
     layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iftrue;
     layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_return_output := layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_return_output;

     -- layer2_node9_MUX[bit_math_h_l1185_c3_9e4b] LATENCY=0
     -- Inputs
     layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_cond <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_cond;
     layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iftrue <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iftrue;
     layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iffalse <= VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_iffalse;
     -- Outputs
     VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_return_output := layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_return_output;

     -- layer2_node1_MUX[bit_math_h_l1097_c3_1a30] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l1097_c3_1a30_cond <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_cond;
     layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iftrue;
     layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_return_output := layer2_node1_MUX_bit_math_h_l1097_c3_1a30_return_output;

     -- layer2_node4_MUX[bit_math_h_l1130_c3_7e5b] LATENCY=0
     -- Inputs
     layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_cond <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_cond;
     layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iftrue <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iftrue;
     layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iffalse <= VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_iffalse;
     -- Outputs
     VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_return_output := layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_return_output;

     -- layer2_node12_MUX[bit_math_h_l1218_c3_fc60] LATENCY=0
     -- Inputs
     layer2_node12_MUX_bit_math_h_l1218_c3_fc60_cond <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_cond;
     layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iftrue <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iftrue;
     layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iffalse <= VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_iffalse;
     -- Outputs
     VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_return_output := layer2_node12_MUX_bit_math_h_l1218_c3_fc60_return_output;

     -- layer2_node15_MUX[bit_math_h_l1251_c3_ecd2] LATENCY=0
     -- Inputs
     layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_cond <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_cond;
     layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iftrue <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iftrue;
     layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iffalse <= VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_iffalse;
     -- Outputs
     VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_return_output := layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_return_output;

     -- layer2_node5_MUX[bit_math_h_l1141_c3_25de] LATENCY=0
     -- Inputs
     layer2_node5_MUX_bit_math_h_l1141_c3_25de_cond <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_cond;
     layer2_node5_MUX_bit_math_h_l1141_c3_25de_iftrue <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_iftrue;
     layer2_node5_MUX_bit_math_h_l1141_c3_25de_iffalse <= VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_iffalse;
     -- Outputs
     VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_return_output := layer2_node5_MUX_bit_math_h_l1141_c3_25de_return_output;

     -- layer2_node10_MUX[bit_math_h_l1196_c3_3974] LATENCY=0
     -- Inputs
     layer2_node10_MUX_bit_math_h_l1196_c3_3974_cond <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_cond;
     layer2_node10_MUX_bit_math_h_l1196_c3_3974_iftrue <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_iftrue;
     layer2_node10_MUX_bit_math_h_l1196_c3_3974_iffalse <= VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_iffalse;
     -- Outputs
     VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_return_output := layer2_node10_MUX_bit_math_h_l1196_c3_3974_return_output;

     -- layer2_node14_MUX[bit_math_h_l1240_c3_75b9] LATENCY=0
     -- Inputs
     layer2_node14_MUX_bit_math_h_l1240_c3_75b9_cond <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_cond;
     layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iftrue <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iftrue;
     layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iffalse <= VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_iffalse;
     -- Outputs
     VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_return_output := layer2_node14_MUX_bit_math_h_l1240_c3_75b9_return_output;

     -- layer2_node7_MUX[bit_math_h_l1163_c3_9403] LATENCY=0
     -- Inputs
     layer2_node7_MUX_bit_math_h_l1163_c3_9403_cond <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_cond;
     layer2_node7_MUX_bit_math_h_l1163_c3_9403_iftrue <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_iftrue;
     layer2_node7_MUX_bit_math_h_l1163_c3_9403_iffalse <= VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_iffalse;
     -- Outputs
     VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_return_output := layer2_node7_MUX_bit_math_h_l1163_c3_9403_return_output;

     -- layer2_node13_MUX[bit_math_h_l1229_c3_6c25] LATENCY=0
     -- Inputs
     layer2_node13_MUX_bit_math_h_l1229_c3_6c25_cond <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_cond;
     layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iftrue <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iftrue;
     layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iffalse <= VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_iffalse;
     -- Outputs
     VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_return_output := layer2_node13_MUX_bit_math_h_l1229_c3_6c25_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_iffalse := VAR_layer2_node0_MUX_bit_math_h_l1086_c3_f1d8_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iffalse := VAR_layer2_node10_MUX_bit_math_h_l1196_c3_3974_return_output;
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iftrue := VAR_layer2_node11_MUX_bit_math_h_l1207_c3_80d7_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_iffalse := VAR_layer2_node12_MUX_bit_math_h_l1218_c3_fc60_return_output;
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_iftrue := VAR_layer2_node13_MUX_bit_math_h_l1229_c3_6c25_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iffalse := VAR_layer2_node14_MUX_bit_math_h_l1240_c3_75b9_return_output;
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iftrue := VAR_layer2_node15_MUX_bit_math_h_l1251_c3_ecd2_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_iftrue := VAR_layer2_node1_MUX_bit_math_h_l1097_c3_1a30_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iffalse := VAR_layer2_node2_MUX_bit_math_h_l1108_c3_0b56_return_output;
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iftrue := VAR_layer2_node3_MUX_bit_math_h_l1119_c3_7df6_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iffalse := VAR_layer2_node4_MUX_bit_math_h_l1130_c3_7e5b_return_output;
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iftrue := VAR_layer2_node5_MUX_bit_math_h_l1141_c3_25de_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iffalse := VAR_layer2_node6_MUX_bit_math_h_l1152_c3_be62_return_output;
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iftrue := VAR_layer2_node7_MUX_bit_math_h_l1163_c3_9403_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iffalse := VAR_layer2_node8_MUX_bit_math_h_l1174_c3_918c_return_output;
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iftrue := VAR_layer2_node9_MUX_bit_math_h_l1185_c3_9e4b_return_output;
     -- layer3_node6_MUX[bit_math_h_l1334_c3_483e] LATENCY=0
     -- Inputs
     layer3_node6_MUX_bit_math_h_l1334_c3_483e_cond <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_cond;
     layer3_node6_MUX_bit_math_h_l1334_c3_483e_iftrue <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_iftrue;
     layer3_node6_MUX_bit_math_h_l1334_c3_483e_iffalse <= VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_iffalse;
     -- Outputs
     VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_return_output := layer3_node6_MUX_bit_math_h_l1334_c3_483e_return_output;

     -- layer3_node2_MUX[bit_math_h_l1290_c3_c56d] LATENCY=0
     -- Inputs
     layer3_node2_MUX_bit_math_h_l1290_c3_c56d_cond <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_cond;
     layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iftrue <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iftrue;
     layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iffalse <= VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_iffalse;
     -- Outputs
     VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_return_output := layer3_node2_MUX_bit_math_h_l1290_c3_c56d_return_output;

     -- layer3_node5_MUX[bit_math_h_l1323_c3_75a2] LATENCY=0
     -- Inputs
     layer3_node5_MUX_bit_math_h_l1323_c3_75a2_cond <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_cond;
     layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iftrue <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iftrue;
     layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iffalse <= VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_iffalse;
     -- Outputs
     VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_return_output := layer3_node5_MUX_bit_math_h_l1323_c3_75a2_return_output;

     -- layer3_node0_MUX[bit_math_h_l1268_c3_324b] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l1268_c3_324b_cond <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_cond;
     layer3_node0_MUX_bit_math_h_l1268_c3_324b_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_iftrue;
     layer3_node0_MUX_bit_math_h_l1268_c3_324b_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_return_output := layer3_node0_MUX_bit_math_h_l1268_c3_324b_return_output;

     -- layer3_node4_MUX[bit_math_h_l1312_c3_4b99] LATENCY=0
     -- Inputs
     layer3_node4_MUX_bit_math_h_l1312_c3_4b99_cond <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_cond;
     layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iftrue <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iftrue;
     layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iffalse <= VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_iffalse;
     -- Outputs
     VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_return_output := layer3_node4_MUX_bit_math_h_l1312_c3_4b99_return_output;

     -- layer3_node1_MUX[bit_math_h_l1279_c3_eea1] LATENCY=0
     -- Inputs
     layer3_node1_MUX_bit_math_h_l1279_c3_eea1_cond <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_cond;
     layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iftrue <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iftrue;
     layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iffalse <= VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_iffalse;
     -- Outputs
     VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_return_output := layer3_node1_MUX_bit_math_h_l1279_c3_eea1_return_output;

     -- layer3_node7_MUX[bit_math_h_l1345_c3_7c85] LATENCY=0
     -- Inputs
     layer3_node7_MUX_bit_math_h_l1345_c3_7c85_cond <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_cond;
     layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iftrue <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iftrue;
     layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iffalse <= VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_iffalse;
     -- Outputs
     VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_return_output := layer3_node7_MUX_bit_math_h_l1345_c3_7c85_return_output;

     -- layer3_node3_MUX[bit_math_h_l1301_c3_98b1] LATENCY=0
     -- Inputs
     layer3_node3_MUX_bit_math_h_l1301_c3_98b1_cond <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_cond;
     layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iftrue <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iftrue;
     layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iffalse <= VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_iffalse;
     -- Outputs
     VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_return_output := layer3_node3_MUX_bit_math_h_l1301_c3_98b1_return_output;

     -- Submodule level 5
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iffalse := VAR_layer3_node0_MUX_bit_math_h_l1268_c3_324b_return_output;
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iftrue := VAR_layer3_node1_MUX_bit_math_h_l1279_c3_eea1_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_iffalse := VAR_layer3_node2_MUX_bit_math_h_l1290_c3_c56d_return_output;
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_iftrue := VAR_layer3_node3_MUX_bit_math_h_l1301_c3_98b1_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_iffalse := VAR_layer3_node4_MUX_bit_math_h_l1312_c3_4b99_return_output;
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_iftrue := VAR_layer3_node5_MUX_bit_math_h_l1323_c3_75a2_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iffalse := VAR_layer3_node6_MUX_bit_math_h_l1334_c3_483e_return_output;
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iftrue := VAR_layer3_node7_MUX_bit_math_h_l1345_c3_7c85_return_output;
     -- layer4_node0_MUX[bit_math_h_l1362_c3_bbba] LATENCY=0
     -- Inputs
     layer4_node0_MUX_bit_math_h_l1362_c3_bbba_cond <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_cond;
     layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iftrue <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iftrue;
     layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iffalse <= VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_iffalse;
     -- Outputs
     VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_return_output := layer4_node0_MUX_bit_math_h_l1362_c3_bbba_return_output;

     -- layer4_node1_MUX[bit_math_h_l1373_c3_31df] LATENCY=0
     -- Inputs
     layer4_node1_MUX_bit_math_h_l1373_c3_31df_cond <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_cond;
     layer4_node1_MUX_bit_math_h_l1373_c3_31df_iftrue <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_iftrue;
     layer4_node1_MUX_bit_math_h_l1373_c3_31df_iffalse <= VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_iffalse;
     -- Outputs
     VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_return_output := layer4_node1_MUX_bit_math_h_l1373_c3_31df_return_output;

     -- layer4_node3_MUX[bit_math_h_l1395_c3_fa88] LATENCY=0
     -- Inputs
     layer4_node3_MUX_bit_math_h_l1395_c3_fa88_cond <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_cond;
     layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iftrue <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iftrue;
     layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iffalse <= VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_iffalse;
     -- Outputs
     VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_return_output := layer4_node3_MUX_bit_math_h_l1395_c3_fa88_return_output;

     -- layer4_node2_MUX[bit_math_h_l1384_c3_d801] LATENCY=0
     -- Inputs
     layer4_node2_MUX_bit_math_h_l1384_c3_d801_cond <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_cond;
     layer4_node2_MUX_bit_math_h_l1384_c3_d801_iftrue <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_iftrue;
     layer4_node2_MUX_bit_math_h_l1384_c3_d801_iffalse <= VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_iffalse;
     -- Outputs
     VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_return_output := layer4_node2_MUX_bit_math_h_l1384_c3_d801_return_output;

     -- Submodule level 6
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iffalse := VAR_layer4_node0_MUX_bit_math_h_l1362_c3_bbba_return_output;
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iftrue := VAR_layer4_node1_MUX_bit_math_h_l1373_c3_31df_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iffalse := VAR_layer4_node2_MUX_bit_math_h_l1384_c3_d801_return_output;
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iftrue := VAR_layer4_node3_MUX_bit_math_h_l1395_c3_fa88_return_output;
     -- layer5_node1_MUX[bit_math_h_l1423_c3_93d3] LATENCY=0
     -- Inputs
     layer5_node1_MUX_bit_math_h_l1423_c3_93d3_cond <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_cond;
     layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iftrue <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iftrue;
     layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iffalse <= VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_iffalse;
     -- Outputs
     VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_return_output := layer5_node1_MUX_bit_math_h_l1423_c3_93d3_return_output;

     -- layer5_node0_MUX[bit_math_h_l1412_c3_ee13] LATENCY=0
     -- Inputs
     layer5_node0_MUX_bit_math_h_l1412_c3_ee13_cond <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_cond;
     layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iftrue <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iftrue;
     layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iffalse <= VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_iffalse;
     -- Outputs
     VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_return_output := layer5_node0_MUX_bit_math_h_l1412_c3_ee13_return_output;

     -- Submodule level 7
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iffalse := VAR_layer5_node0_MUX_bit_math_h_l1412_c3_ee13_return_output;
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iftrue := VAR_layer5_node1_MUX_bit_math_h_l1423_c3_93d3_return_output;
     -- layer6_node0_MUX[bit_math_h_l1440_c3_08eb] LATENCY=0
     -- Inputs
     layer6_node0_MUX_bit_math_h_l1440_c3_08eb_cond <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_cond;
     layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iftrue <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iftrue;
     layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iffalse <= VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_iffalse;
     -- Outputs
     VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_return_output := layer6_node0_MUX_bit_math_h_l1440_c3_08eb_return_output;

     -- Submodule level 8
     VAR_return_output := VAR_layer6_node0_MUX_bit_math_h_l1440_c3_08eb_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
