-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2640_c6_d665]
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2640_c2_58df]
signal n8_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2640_c2_58df]
signal t8_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2640_c2_58df]
signal l8_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2640_c2_58df]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2653_c11_7ebb]
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2653_c7_2a26]
signal n8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2653_c7_2a26]
signal t8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2653_c7_2a26]
signal l8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2653_c7_2a26]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2653_c7_2a26]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2653_c7_2a26]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2653_c7_2a26]
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2653_c7_2a26]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2656_c11_1348]
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2656_c7_deee]
signal n8_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2656_c7_deee]
signal t8_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2656_c7_deee]
signal l8_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c7_deee]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c7_deee]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c7_deee]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2656_c7_deee]
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c7_deee]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2660_c11_a4bb]
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2660_c7_8db8]
signal n8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(7 downto 0);

-- l8_MUX[uxn_opcodes_h_l2660_c7_8db8]
signal l8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2660_c7_8db8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2660_c7_8db8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2660_c7_8db8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2660_c7_8db8]
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2660_c7_8db8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2662_c30_9b4e]
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2667_c11_c401]
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2667_c7_6f7f]
signal l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2667_c7_6f7f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2667_c7_6f7f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2667_c7_6f7f]
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2667_c7_6f7f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_5c28]
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_ca51]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_ca51]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_ca51]
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a6df( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_ram_write := ref_toks_8;
      base.is_stack_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_left,
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_right,
BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output);

-- n8_MUX_uxn_opcodes_h_l2640_c2_58df
n8_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
n8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
n8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
n8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- t8_MUX_uxn_opcodes_h_l2640_c2_58df
t8_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
t8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
t8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
t8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- l8_MUX_uxn_opcodes_h_l2640_c2_58df
l8_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
l8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
l8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
l8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_left,
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_right,
BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output);

-- n8_MUX_uxn_opcodes_h_l2653_c7_2a26
n8_MUX_uxn_opcodes_h_l2653_c7_2a26 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond,
n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue,
n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse,
n8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output);

-- t8_MUX_uxn_opcodes_h_l2653_c7_2a26
t8_MUX_uxn_opcodes_h_l2653_c7_2a26 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond,
t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue,
t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse,
t8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output);

-- l8_MUX_uxn_opcodes_h_l2653_c7_2a26
l8_MUX_uxn_opcodes_h_l2653_c7_2a26 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond,
l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue,
l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse,
l8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_cond,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_left,
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_right,
BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output);

-- n8_MUX_uxn_opcodes_h_l2656_c7_deee
n8_MUX_uxn_opcodes_h_l2656_c7_deee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2656_c7_deee_cond,
n8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue,
n8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse,
n8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output);

-- t8_MUX_uxn_opcodes_h_l2656_c7_deee
t8_MUX_uxn_opcodes_h_l2656_c7_deee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2656_c7_deee_cond,
t8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue,
t8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse,
t8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output);

-- l8_MUX_uxn_opcodes_h_l2656_c7_deee
l8_MUX_uxn_opcodes_h_l2656_c7_deee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2656_c7_deee_cond,
l8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue,
l8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse,
l8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_cond,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_left,
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_right,
BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output);

-- n8_MUX_uxn_opcodes_h_l2660_c7_8db8
n8_MUX_uxn_opcodes_h_l2660_c7_8db8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond,
n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue,
n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse,
n8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output);

-- l8_MUX_uxn_opcodes_h_l2660_c7_8db8
l8_MUX_uxn_opcodes_h_l2660_c7_8db8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond,
l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue,
l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse,
l8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e
sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_ins,
sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_x,
sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_y,
sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_left,
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_right,
BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output);

-- l8_MUX_uxn_opcodes_h_l2667_c7_6f7f
l8_MUX_uxn_opcodes_h_l2667_c7_6f7f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond,
l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue,
l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse,
l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_left,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_right,
BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_cond,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output,
 n8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 t8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 l8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output,
 n8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output,
 t8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output,
 l8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output,
 n8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output,
 t8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output,
 l8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output,
 n8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output,
 l8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output,
 sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output,
 l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_4529 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_6017 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_504d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_b37b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_654b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_f955 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_0358 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_178c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_ca51_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_6408_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_441e_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2656_l2653_l2673_l2667_l2660_DUPLICATE_8623_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2653_l2656_l2660_DUPLICATE_43bb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2636_l2679_DUPLICATE_27b0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_654b := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2664_c3_654b;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_4529 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2645_c3_4529;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_right := to_unsigned(2, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_178c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2674_c3_178c;
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_504d := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2654_c3_504d;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_6017 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2650_c3_6017;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_b37b := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2657_c3_b37b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_f955 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2669_c3_f955;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_0358 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_0358;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse := t8;
     -- sp_relative_shift[uxn_opcodes_h_l2662_c30_9b4e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_ins;
     sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_x;
     sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_return_output := sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2656_c11_1348] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_left;
     BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output := BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_441e LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_441e_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2640_c6_d665] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_left;
     BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output := BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_6408 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_6408_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2653_l2656_l2660_DUPLICATE_43bb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2653_l2656_l2660_DUPLICATE_43bb_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2673_c11_5c28] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_left;
     BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output := BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2653_c11_7ebb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2673_c7_ca51] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_ca51_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2656_l2653_l2673_l2667_l2660_DUPLICATE_8623 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2656_l2653_l2673_l2667_l2660_DUPLICATE_8623_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2660_c11_a4bb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_left;
     BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output := BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2667_c11_c401] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_left;
     BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output := BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_58df_return_output := result.is_stack_index_flipped;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_58df_return_output := result.is_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_58df_return_output := result.is_vram_write;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_58df_return_output := result.is_pc_updated;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2640_c6_d665_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2653_c11_7ebb_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c11_1348_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2660_c11_a4bb_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2667_c11_c401_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2673_c11_5c28_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_441e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_441e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2653_l2667_l2656_DUPLICATE_441e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2656_l2653_l2673_l2667_l2660_DUPLICATE_8623_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2656_l2653_l2673_l2667_l2660_DUPLICATE_8623_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2656_l2653_l2673_l2667_l2660_DUPLICATE_8623_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2656_l2653_l2673_l2667_l2660_DUPLICATE_8623_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2656_l2653_l2673_l2667_l2660_DUPLICATE_8623_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2653_l2656_l2660_DUPLICATE_43bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2653_l2656_l2660_DUPLICATE_43bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2653_l2656_l2660_DUPLICATE_43bb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_6408_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_6408_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_6408_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2653_l2656_l2673_l2640_DUPLICATE_6408_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2640_c2_58df_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2640_c2_58df_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2640_c2_58df_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2640_c2_58df_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2673_c7_ca51_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2662_c30_9b4e_return_output;
     -- n8_MUX[uxn_opcodes_h_l2660_c7_8db8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond;
     n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue;
     n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output := n8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2673_c7_ca51] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output := result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output;

     -- l8_MUX[uxn_opcodes_h_l2667_c7_6f7f] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond;
     l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue;
     l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output := l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2673_c7_ca51] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2667_c7_6f7f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- t8_MUX[uxn_opcodes_h_l2656_c7_deee] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2656_c7_deee_cond <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_cond;
     t8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue;
     t8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output := t8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2673_c7_ca51] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2660_c7_8db8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2673_c7_ca51_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;
     -- l8_MUX[uxn_opcodes_h_l2660_c7_8db8] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_cond;
     l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue;
     l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output := l8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2667_c7_6f7f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2660_c7_8db8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2667_c7_6f7f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2667_c7_6f7f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;

     -- n8_MUX[uxn_opcodes_h_l2656_c7_deee] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2656_c7_deee_cond <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_cond;
     n8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue;
     n8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output := n8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;

     -- t8_MUX[uxn_opcodes_h_l2653_c7_2a26] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond;
     t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue;
     t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output := t8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c7_deee] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2667_c7_6f7f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c7_deee] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2660_c7_8db8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;

     -- t8_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     t8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     t8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := t8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2653_c7_2a26] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2660_c7_8db8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2653_c7_2a26] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond;
     n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue;
     n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output := n8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;

     -- l8_MUX[uxn_opcodes_h_l2656_c7_deee] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2656_c7_deee_cond <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_cond;
     l8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue;
     l8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output := l8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2660_c7_8db8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2660_c7_8db8_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;
     -- n8_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     n8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     n8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := n8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c7_deee] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c7_deee] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2653_c7_2a26] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;

     -- l8_MUX[uxn_opcodes_h_l2653_c7_2a26] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_cond;
     l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue;
     l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output := l8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2656_c7_deee] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_return_output := result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c7_deee_return_output;
     -- l8_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     l8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     l8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := l8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2653_c7_2a26] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2653_c7_2a26] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output := result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2653_c7_2a26] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2653_c7_2a26_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2640_c2_58df] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2636_l2679_DUPLICATE_27b0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2636_l2679_DUPLICATE_27b0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a6df(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2640_c2_58df_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2636_l2679_DUPLICATE_27b0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a6df_uxn_opcodes_h_l2636_l2679_DUPLICATE_27b0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
