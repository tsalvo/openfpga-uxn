-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 33
entity VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
port(
 elem_val : in unsigned(7 downto 0);
 ref_toks_0 : in uint8_t_16;
 var_dim_0 : in unsigned(3 downto 0);
 return_output : out uint8_t_array_16_t);
end VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28;
architecture arch of VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_0CLK_6481cb28 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_return_output : unsigned(0 downto 0);

-- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105]
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_cond : unsigned(0 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iftrue : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iffalse : unsigned(7 downto 0);
signal rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_return_output : unsigned(0 downto 0);

-- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48]
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_cond : unsigned(0 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iftrue : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iffalse : unsigned(7 downto 0);
signal rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_return_output : unsigned(0 downto 0);

-- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416]
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_cond : unsigned(0 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iftrue : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iffalse : unsigned(7 downto 0);
signal rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_return_output : unsigned(0 downto 0);

-- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd]
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_cond : unsigned(0 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iftrue : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iffalse : unsigned(7 downto 0);
signal rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_return_output : unsigned(0 downto 0);

-- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b]
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_cond : unsigned(0 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iftrue : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iffalse : unsigned(7 downto 0);
signal rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_return_output : unsigned(0 downto 0);

-- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53]
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_cond : unsigned(0 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iftrue : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iffalse : unsigned(7 downto 0);
signal rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_return_output : unsigned(0 downto 0);

-- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8]
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_cond : unsigned(0 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iftrue : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iffalse : unsigned(7 downto 0);
signal rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_return_output : unsigned(0 downto 0);

-- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5]
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_cond : unsigned(0 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iftrue : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iffalse : unsigned(7 downto 0);
signal rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_right : unsigned(1 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_return_output : unsigned(0 downto 0);

-- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf]
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_cond : unsigned(0 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iftrue : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iffalse : unsigned(7 downto 0);
signal rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_return_output : unsigned(0 downto 0);

-- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141]
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_cond : unsigned(0 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iftrue : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iffalse : unsigned(7 downto 0);
signal rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_return_output : unsigned(0 downto 0);

-- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09]
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_cond : unsigned(0 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iftrue : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iffalse : unsigned(7 downto 0);
signal rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_return_output : unsigned(0 downto 0);

-- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90]
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_cond : unsigned(0 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iftrue : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iffalse : unsigned(7 downto 0);
signal rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_return_output : unsigned(0 downto 0);

-- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287]
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_cond : unsigned(0 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iftrue : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iffalse : unsigned(7 downto 0);
signal rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_right : unsigned(0 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_return_output : unsigned(0 downto 0);

-- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27]
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_cond : unsigned(0 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iftrue : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iffalse : unsigned(7 downto 0);
signal rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_right : unsigned(2 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_return_output : unsigned(0 downto 0);

-- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf]
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_cond : unsigned(0 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iftrue : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iffalse : unsigned(7 downto 0);
signal rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28]
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_left : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_right : unsigned(3 downto 0);
signal BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_return_output : unsigned(0 downto 0);

-- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b]
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_cond : unsigned(0 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iftrue : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iffalse : unsigned(7 downto 0);
signal rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_return_output : unsigned(7 downto 0);

function CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_80e1( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_array_16_t is
 
  variable base : uint8_t_array_16_t; 
  variable return_output : uint8_t_array_16_t;
begin
      base.data(10) := ref_toks_0;
      base.data(2) := ref_toks_1;
      base.data(5) := ref_toks_2;
      base.data(11) := ref_toks_3;
      base.data(8) := ref_toks_4;
      base.data(14) := ref_toks_5;
      base.data(0) := ref_toks_6;
      base.data(6) := ref_toks_7;
      base.data(3) := ref_toks_8;
      base.data(9) := ref_toks_9;
      base.data(12) := ref_toks_10;
      base.data(15) := ref_toks_11;
      base.data(4) := ref_toks_12;
      base.data(1) := ref_toks_13;
      base.data(7) := ref_toks_14;
      base.data(13) := ref_toks_15;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_return_output);

-- rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_cond,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iftrue,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iffalse,
rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_return_output);

-- rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_cond,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iftrue,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iffalse,
rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_return_output);

-- rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_cond,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iftrue,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iffalse,
rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_return_output);

-- rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_cond,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iftrue,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iffalse,
rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_return_output);

-- rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_cond,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iftrue,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iffalse,
rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_return_output);

-- rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_cond,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iftrue,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iffalse,
rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_return_output);

-- rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_cond,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iftrue,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iffalse,
rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_return_output);

-- rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_cond,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iftrue,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iffalse,
rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_return_output);

-- rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_cond,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iftrue,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iffalse,
rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_return_output);

-- rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_cond,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iftrue,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iffalse,
rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_return_output);

-- rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_cond,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iftrue,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iffalse,
rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_return_output);

-- rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_cond,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iftrue,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iffalse,
rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_return_output);

-- rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_cond,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iftrue,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iffalse,
rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40 : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_return_output);

-- rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_cond,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iftrue,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iffalse,
rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_return_output);

-- rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_cond,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iftrue,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iffalse,
rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_return_output);

-- BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28 : entity work.BIN_OP_EQ_uint4_t_uint4_t_0CLK_de264c78 port map (
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_left,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_right,
BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_return_output);

-- rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_cond,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iftrue,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iffalse,
rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 elem_val,
 ref_toks_0,
 var_dim_0,
 -- All submodule outputs
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_return_output,
 rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_return_output,
 rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_return_output,
 rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_return_output,
 rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_return_output,
 rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_return_output,
 rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_return_output,
 rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_return_output,
 rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_return_output,
 rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_return_output,
 rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_return_output,
 rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_return_output,
 rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_return_output,
 rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_return_output,
 rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_return_output,
 rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_return_output,
 BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_return_output,
 rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_elem_val : unsigned(7 downto 0);
 variable VAR_ref_toks_0 : uint8_t_16;
 variable VAR_var_dim_0 : unsigned(3 downto 0);
 variable VAR_return_output : uint8_t_array_16_t;
 variable VAR_base : uint8_t_16;
 variable VAR_rv : uint8_t_array_16_t;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c16_3140_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_5f08_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_c21d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_9c2d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c15_203c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c16_bac0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_fb22_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_e5d6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_b1fb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c15_3871_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_76b4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c16_d1c7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_8ee9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_4d1e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c15_0c2f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_f81e_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_right : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_return_output : unsigned(0 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iftrue : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iffalse : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_return_output : unsigned(7 downto 0);
 variable VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_80e1_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_4e84_return_output : uint8_t_array_16_t;
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_right := to_unsigned(10, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_right := to_unsigned(13, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_right := to_unsigned(6, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_right := to_unsigned(15, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_right := to_unsigned(11, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_right := to_unsigned(8, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_right := to_unsigned(12, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_right := to_unsigned(7, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_right := to_unsigned(9, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_right := to_unsigned(14, 4);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_right := to_unsigned(3, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_elem_val := elem_val;
     VAR_ref_toks_0 := ref_toks_0;
     VAR_var_dim_0 := var_dim_0;

     -- Submodule level 0
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iftrue := VAR_elem_val;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iftrue := VAR_elem_val;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iftrue := VAR_elem_val;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iftrue := VAR_elem_val;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iftrue := VAR_elem_val;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iftrue := VAR_elem_val;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iftrue := VAR_elem_val;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iftrue := VAR_elem_val;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iftrue := VAR_elem_val;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iftrue := VAR_elem_val;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iftrue := VAR_elem_val;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iftrue := VAR_elem_val;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iftrue := VAR_elem_val;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iftrue := VAR_elem_val;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iftrue := VAR_elem_val;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iftrue := VAR_elem_val;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_left := VAR_var_dim_0;
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_left := VAR_var_dim_0;
     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_3_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_b1fb] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_b1fb_return_output := VAR_ref_toks_0(3);

     -- CONST_REF_RD_uint8_t_uint8_t_16_4_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_8ee9] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_8ee9_return_output := VAR_ref_toks_0(4);

     -- CONST_REF_RD_uint8_t_uint8_t_16_1_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_4d1e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_4d1e_return_output := VAR_ref_toks_0(1);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_10_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c16_3140] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c16_3140_return_output := VAR_ref_toks_0(10);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_11_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_9c2d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_9c2d_return_output := VAR_ref_toks_0(11);

     -- CONST_REF_RD_uint8_t_uint8_t_16_13_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_f81e] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_f81e_return_output := VAR_ref_toks_0(13);

     -- CONST_REF_RD_uint8_t_uint8_t_16_12_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_76b4] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_76b4_return_output := VAR_ref_toks_0(12);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_6_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_e5d6] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_e5d6_return_output := VAR_ref_toks_0(6);

     -- CONST_REF_RD_uint8_t_uint8_t_16_0_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_fb22] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_fb22_return_output := VAR_ref_toks_0(0);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_5_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_c21d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_c21d_return_output := VAR_ref_toks_0(5);

     -- CONST_REF_RD_uint8_t_uint8_t_16_14_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c16_bac0] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c16_bac0_return_output := VAR_ref_toks_0(14);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_return_output;

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_8_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c15_203c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c15_203c_return_output := VAR_ref_toks_0(8);

     -- CONST_REF_RD_uint8_t_uint8_t_16_15_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c16_d1c7] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c16_d1c7_return_output := VAR_ref_toks_0(15);

     -- CONST_REF_RD_uint8_t_uint8_t_16_2_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_5f08] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_5f08_return_output := VAR_ref_toks_0(2);

     -- CONST_REF_RD_uint8_t_uint8_t_16_7_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c15_0c2f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c15_0c2f_return_output := VAR_ref_toks_0(7);

     -- BIN_OP_EQ[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465] LATENCY=0
     -- Inputs
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_left <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_left;
     BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_right <= VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_right;
     -- Outputs
     VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_return_output := BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_16_9_d41d[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c15_3871] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c15_3871_return_output := VAR_ref_toks_0(9);

     -- Submodule level 1
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l105_c5_f811_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l111_c5_be40_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l117_c5_f465_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l123_c5_3c28_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l33_c5_4bb5_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l39_c5_f08c_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l45_c5_d824_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l51_c5_e64b_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l57_c5_afc2_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l63_c5_7f13_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l69_c5_17de_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l75_c5_0ce5_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l81_c5_8e64_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l87_c5_10ce_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l93_c5_618f_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_cond := VAR_BIN_OP_EQ_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l99_c5_18ce_return_output;
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_0_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l21_c15_fb22_return_output;
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_10_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l15_c16_3140_return_output;
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_11_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l18_c16_9c2d_return_output;
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_12_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l25_c16_76b4_return_output;
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_13_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l30_c16_f81e_return_output;
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_14_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l20_c16_bac0_return_output;
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_15_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l26_c16_d1c7_return_output;
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_1_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l28_c15_4d1e_return_output;
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_2_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l16_c15_5f08_return_output;
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_3_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l23_c15_b1fb_return_output;
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_4_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l27_c15_8ee9_return_output;
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_5_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l17_c15_c21d_return_output;
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_6_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l22_c15_e5d6_return_output;
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_7_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l29_c15_0c2f_return_output;
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_8_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l19_c15_203c_return_output;
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_16_9_d41d_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l24_c15_3871_return_output;
     -- rv_data_4_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287] LATENCY=0
     -- Inputs
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_cond <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_cond;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iftrue <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iftrue;
     rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iffalse <= VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_iffalse;
     -- Outputs
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_return_output := rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_return_output;

     -- rv_data_5_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416] LATENCY=0
     -- Inputs
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_cond <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_cond;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iftrue <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iftrue;
     rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iffalse <= VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_iffalse;
     -- Outputs
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_return_output := rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_return_output;

     -- rv_data_6_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5] LATENCY=0
     -- Inputs
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_cond <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_cond;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iftrue <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iftrue;
     rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iffalse <= VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_iffalse;
     -- Outputs
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_return_output := rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_return_output;

     -- rv_data_15_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90] LATENCY=0
     -- Inputs
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_cond <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_cond;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iftrue <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iftrue;
     rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iffalse <= VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_iffalse;
     -- Outputs
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_return_output := rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_return_output;

     -- rv_data_12_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09] LATENCY=0
     -- Inputs
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_cond <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_cond;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iftrue <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iftrue;
     rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iffalse <= VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_iffalse;
     -- Outputs
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_return_output := rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_return_output;

     -- rv_data_0_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8] LATENCY=0
     -- Inputs
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_cond <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_cond;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iftrue <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iftrue;
     rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iffalse <= VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_iffalse;
     -- Outputs
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_return_output := rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_return_output;

     -- rv_data_7_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf] LATENCY=0
     -- Inputs
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_cond <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_cond;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iftrue <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iftrue;
     rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iffalse <= VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_iffalse;
     -- Outputs
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_return_output := rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_return_output;

     -- rv_data_3_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf] LATENCY=0
     -- Inputs
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_cond <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_cond;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iftrue <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iftrue;
     rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iffalse <= VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_iffalse;
     -- Outputs
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_return_output := rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_return_output;

     -- rv_data_11_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd] LATENCY=0
     -- Inputs
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_cond <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_cond;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iftrue <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iftrue;
     rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iffalse <= VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_iffalse;
     -- Outputs
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_return_output := rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_return_output;

     -- rv_data_9_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141] LATENCY=0
     -- Inputs
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_cond <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_cond;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iftrue <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iftrue;
     rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iffalse <= VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_iffalse;
     -- Outputs
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_return_output := rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_return_output;

     -- rv_data_1_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27] LATENCY=0
     -- Inputs
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_cond <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_cond;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iftrue <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iftrue;
     rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iffalse <= VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_iffalse;
     -- Outputs
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_return_output := rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_return_output;

     -- rv_data_14_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53] LATENCY=0
     -- Inputs
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_cond <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_cond;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iftrue <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iftrue;
     rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iffalse <= VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_iffalse;
     -- Outputs
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_return_output := rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_return_output;

     -- rv_data_13_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b] LATENCY=0
     -- Inputs
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_cond <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_cond;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iftrue <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iftrue;
     rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iffalse <= VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_iffalse;
     -- Outputs
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_return_output := rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_return_output;

     -- rv_data_10_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105] LATENCY=0
     -- Inputs
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_cond <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_cond;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iftrue <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iftrue;
     rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iffalse <= VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_iffalse;
     -- Outputs
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_return_output := rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_return_output;

     -- rv_data_8_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b] LATENCY=0
     -- Inputs
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_cond <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_cond;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iftrue <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iftrue;
     rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iffalse <= VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_iffalse;
     -- Outputs
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_return_output := rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_return_output;

     -- rv_data_2_MUX[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48] LATENCY=0
     -- Inputs
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_cond <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_cond;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iftrue <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iftrue;
     rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iffalse <= VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_iffalse;
     -- Outputs
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_return_output := rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_return_output;

     -- Submodule level 2
     -- CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_80e1[VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_4e84] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_80e1_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_4e84_return_output := CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_80e1(
     VAR_rv_data_10_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l32_c2_7105_return_output,
     VAR_rv_data_2_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l38_c2_4d48_return_output,
     VAR_rv_data_5_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l44_c2_7416_return_output,
     VAR_rv_data_11_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l50_c2_b4fd_return_output,
     VAR_rv_data_8_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l56_c2_e34b_return_output,
     VAR_rv_data_14_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l62_c2_dd53_return_output,
     VAR_rv_data_0_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l68_c2_8bd8_return_output,
     VAR_rv_data_6_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l74_c2_97b5_return_output,
     VAR_rv_data_3_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l80_c2_7fdf_return_output,
     VAR_rv_data_9_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l86_c2_0141_return_output,
     VAR_rv_data_12_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l92_c2_bb09_return_output,
     VAR_rv_data_15_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l98_c2_6b90_return_output,
     VAR_rv_data_4_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l104_c2_f287_return_output,
     VAR_rv_data_1_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l110_c2_6c27_return_output,
     VAR_rv_data_7_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l116_c2_3caf_return_output,
     VAR_rv_data_13_MUX_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l122_c2_057b_return_output);

     -- Submodule level 3
     VAR_return_output := VAR_CONST_REF_RD_uint8_t_array_16_t_uint8_t_array_16_t_80e1_VAR_REF_ASSIGN_uint8_t_uint8_t_16_VAR_7a60_c_l129_c10_4e84_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
