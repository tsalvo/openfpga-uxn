-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity nip2_0CLK_9a874500 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end nip2_0CLK_9a874500;
architecture arch of nip2_0CLK_9a874500 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2061_c6_d790]
signal BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2061_c1_1ccc]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2061_c2_01c0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2061_c2_01c0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2061_c2_01c0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2061_c2_01c0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2061_c2_01c0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2061_c2_01c0]
signal result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2061_c2_01c0]
signal t16_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(15 downto 0);

-- printf_uxn_opcodes_h_l2062_c3_0425[uxn_opcodes_h_l2062_c3_0425]
signal printf_uxn_opcodes_h_l2062_c3_0425_uxn_opcodes_h_l2062_c3_0425_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2066_c11_b250]
signal BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2066_c7_4924]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2066_c7_4924]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2066_c7_4924]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2066_c7_4924]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2066_c7_4924]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2066_c7_4924]
signal result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2066_c7_4924]
signal t16_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2069_c11_a2b0]
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2069_c7_3bd8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2069_c7_3bd8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2069_c7_3bd8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2069_c7_3bd8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2069_c7_3bd8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2069_c7_3bd8]
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2069_c7_3bd8]
signal t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2071_c3_b9e4]
signal CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2073_c11_e3b0]
signal BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2073_c7_9aed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2073_c7_9aed]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2073_c7_9aed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2073_c7_9aed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2073_c7_9aed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2073_c7_9aed]
signal result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2073_c7_9aed]
signal t16_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2074_c3_20ce]
signal BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2076_c30_8040]
signal sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2081_c11_ae6c]
signal BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2081_c7_fe24]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2081_c7_fe24]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2081_c7_fe24]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2081_c7_fe24]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2081_c7_fe24]
signal result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(7 downto 0);

-- CONST_SR_8[uxn_opcodes_h_l2084_c31_dad1]
signal CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_x : unsigned(15 downto 0);
signal CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2086_c11_6798]
signal BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2086_c7_c53f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2086_c7_c53f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_8c29( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790
BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_left,
BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_right,
BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0
result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output);

-- t16_MUX_uxn_opcodes_h_l2061_c2_01c0
t16_MUX_uxn_opcodes_h_l2061_c2_01c0 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2061_c2_01c0_cond,
t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue,
t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse,
t16_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output);

-- printf_uxn_opcodes_h_l2062_c3_0425_uxn_opcodes_h_l2062_c3_0425
printf_uxn_opcodes_h_l2062_c3_0425_uxn_opcodes_h_l2062_c3_0425 : entity work.printf_uxn_opcodes_h_l2062_c3_0425_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2062_c3_0425_uxn_opcodes_h_l2062_c3_0425_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250
BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_left,
BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_right,
BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924
result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924
result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924
result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924
result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924
result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_cond,
result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_return_output);

-- t16_MUX_uxn_opcodes_h_l2066_c7_4924
t16_MUX_uxn_opcodes_h_l2066_c7_4924 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2066_c7_4924_cond,
t16_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue,
t16_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse,
t16_MUX_uxn_opcodes_h_l2066_c7_4924_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_left,
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_right,
BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8
result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output);

-- t16_MUX_uxn_opcodes_h_l2069_c7_3bd8
t16_MUX_uxn_opcodes_h_l2069_c7_3bd8 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond,
t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue,
t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse,
t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4
CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_x,
CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0
BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_left,
BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_right,
BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed
result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_cond,
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output);

-- t16_MUX_uxn_opcodes_h_l2073_c7_9aed
t16_MUX_uxn_opcodes_h_l2073_c7_9aed : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2073_c7_9aed_cond,
t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue,
t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse,
t16_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce
BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_left,
BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_right,
BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2076_c30_8040
sp_relative_shift_uxn_opcodes_h_l2076_c30_8040 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_ins,
sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_x,
sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_y,
sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c
BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_left,
BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_right,
BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24
result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24
result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24
result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24
result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_cond,
result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output);

-- CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1
CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1 : entity work.CONST_SR_8_uint16_t_0CLK_de264c78 port map (
CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_x,
CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798
BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_left,
BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_right,
BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f
result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f
result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
 t16_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_return_output,
 t16_MUX_uxn_opcodes_h_l2066_c7_4924_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output,
 t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output,
 CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output,
 t16_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_return_output,
 sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output,
 CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2063_c3_0643 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2062_c3_0425_uxn_opcodes_h_l2062_c3_0425_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2067_c3_e0cd : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2078_c3_a13c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2079_c21_7b70_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2083_c3_e716 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_cond : unsigned(0 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_x : unsigned(15 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2084_c21_0883_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_40dd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2086_l2081_l2069_l2066_DUPLICATE_855b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2061_l2073_l2066_DUPLICATE_5797_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_ea5e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2086_l2081_l2073_l2069_l2066_DUPLICATE_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2074_l2070_DUPLICATE_1b78_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2069_l2081_DUPLICATE_fa4f_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2057_l2091_DUPLICATE_bc14_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2063_c3_0643 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2063_c3_0643;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_right := to_unsigned(4, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_right := to_unsigned(5, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2067_c3_e0cd := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2067_c3_e0cd;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2078_c3_a13c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2078_c3_a13c;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2083_c3_e716 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2083_c3_e716;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_left := t16;
     VAR_CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_x := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2086_l2081_l2073_l2069_l2066_DUPLICATE_ff6d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2086_l2081_l2073_l2069_l2066_DUPLICATE_ff6d_return_output := result.is_opc_done;

     -- CONST_SR_8[uxn_opcodes_h_l2084_c31_dad1] LATENCY=0
     -- Inputs
     CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_x <= VAR_CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_x;
     -- Outputs
     VAR_CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_return_output := CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2074_l2070_DUPLICATE_1b78 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2074_l2070_DUPLICATE_1b78_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- BIN_OP_EQ[uxn_opcodes_h_l2073_c11_e3b0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2076_c30_8040] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_ins;
     sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_x;
     sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_return_output := sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2081_c11_ae6c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2086_l2081_l2069_l2066_DUPLICATE_855b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2086_l2081_l2069_l2066_DUPLICATE_855b_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_40dd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_40dd_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2061_l2073_l2066_DUPLICATE_5797 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2061_l2073_l2066_DUPLICATE_5797_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2086_c11_6798] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_left;
     BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_return_output := BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2061_c6_d790] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_left;
     BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output := BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_ea5e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_ea5e_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2066_c11_b250] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_left;
     BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output := BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2069_c11_a2b0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2069_l2081_DUPLICATE_fa4f LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2069_l2081_DUPLICATE_fa4f_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2061_c6_d790_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2066_c11_b250_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2069_c11_a2b0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2073_c11_e3b0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2081_c11_ae6c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2086_c11_6798_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2074_l2070_DUPLICATE_1b78_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2074_l2070_DUPLICATE_1b78_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2061_l2073_l2066_DUPLICATE_5797_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2061_l2073_l2066_DUPLICATE_5797_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2061_l2073_l2066_DUPLICATE_5797_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2069_l2061_l2073_l2066_DUPLICATE_5797_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2086_l2081_l2073_l2069_l2066_DUPLICATE_ff6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2086_l2081_l2073_l2069_l2066_DUPLICATE_ff6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2086_l2081_l2073_l2069_l2066_DUPLICATE_ff6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2086_l2081_l2073_l2069_l2066_DUPLICATE_ff6d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2086_l2081_l2073_l2069_l2066_DUPLICATE_ff6d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_40dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_40dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_40dd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_40dd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2086_l2081_l2069_l2066_DUPLICATE_855b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2086_l2081_l2069_l2066_DUPLICATE_855b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2086_l2081_l2069_l2066_DUPLICATE_855b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2086_l2081_l2069_l2066_DUPLICATE_855b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2061_l2086_l2081_l2069_l2066_DUPLICATE_855b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2069_l2081_DUPLICATE_fa4f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2069_l2081_DUPLICATE_fa4f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_ea5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_ea5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_ea5e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2069_l2061_l2066_l2081_DUPLICATE_ea5e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2076_c30_8040_return_output;
     -- CONST_SL_8[uxn_opcodes_h_l2071_c3_b9e4] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_return_output := CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2074_c3_20ce] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_left;
     BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_return_output := BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2084_c21_0883] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2084_c21_0883_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_CONST_SR_8_uxn_opcodes_h_l2084_c31_dad1_return_output);

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2086_c7_c53f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2061_c1_1ccc] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2073_c7_9aed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2081_c7_fe24] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2086_c7_c53f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2081_c7_fe24] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2084_c21_0883_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2071_c3_b9e4_return_output;
     VAR_printf_uxn_opcodes_h_l2062_c3_0425_uxn_opcodes_h_l2062_c3_0425_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2061_c1_1ccc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2086_c7_c53f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2073_c7_9aed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2069_c7_3bd8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2081_c7_fe24] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2081_c7_fe24] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2079_c21_7b70] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2079_c21_7b70_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_BIN_OP_OR_uxn_opcodes_h_l2074_c3_20ce_return_output);

     -- printf_uxn_opcodes_h_l2062_c3_0425[uxn_opcodes_h_l2062_c3_0425] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2062_c3_0425_uxn_opcodes_h_l2062_c3_0425_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2062_c3_0425_uxn_opcodes_h_l2062_c3_0425_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- t16_MUX[uxn_opcodes_h_l2073_c7_9aed] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2073_c7_9aed_cond <= VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_cond;
     t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue;
     t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output := t16_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2073_c7_9aed] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2081_c7_fe24] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output := result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2079_c21_7b70_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2081_c7_fe24_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2069_c7_3bd8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2066_c7_4924] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2069_c7_3bd8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;

     -- t16_MUX[uxn_opcodes_h_l2069_c7_3bd8] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond <= VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond;
     t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue;
     t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output := t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2073_c7_9aed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output := result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2073_c7_9aed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2073_c7_9aed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2073_c7_9aed_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2061_c2_01c0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2069_c7_3bd8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;

     -- t16_MUX[uxn_opcodes_h_l2066_c7_4924] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2066_c7_4924_cond <= VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_cond;
     t16_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue;
     t16_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_return_output := t16_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2069_c7_3bd8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2066_c7_4924] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2069_c7_3bd8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2066_c7_4924] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2069_c7_3bd8_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2061_c2_01c0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2066_c7_4924] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2061_c2_01c0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2066_c7_4924] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2066_c7_4924] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_return_output := result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;

     -- t16_MUX[uxn_opcodes_h_l2061_c2_01c0] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2061_c2_01c0_cond <= VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_cond;
     t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue;
     t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output := t16_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2066_c7_4924_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2061_c2_01c0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2061_c2_01c0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2061_c2_01c0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2057_l2091_DUPLICATE_bc14 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2057_l2091_DUPLICATE_bc14_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_8c29(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2061_c2_01c0_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2057_l2091_DUPLICATE_bc14_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_8c29_uxn_opcodes_h_l2057_l2091_DUPLICATE_bc14_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
