-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity sta_0CLK_bce25fe8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sta_0CLK_bce25fe8;
architecture arch of sta_0CLK_bce25fe8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2316_c6_e0c3]
signal BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(7 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2316_c2_753d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2316_c2_753d]
signal n8_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2316_c2_753d]
signal t16_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2329_c11_75ab]
signal BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2329_c7_cc75]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2329_c7_cc75]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2329_c7_cc75]
signal result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2329_c7_cc75]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2329_c7_cc75]
signal result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2329_c7_cc75]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2329_c7_cc75]
signal n8_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2329_c7_cc75]
signal t16_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2332_c11_93ed]
signal BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2332_c7_2c18]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2332_c7_2c18]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2332_c7_2c18]
signal result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2332_c7_2c18]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2332_c7_2c18]
signal result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2332_c7_2c18]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2332_c7_2c18]
signal n8_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2332_c7_2c18]
signal t16_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l2334_c3_73cc]
signal CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2337_c11_7b3a]
signal BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2337_c7_7acd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2337_c7_7acd]
signal result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2337_c7_7acd]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2337_c7_7acd]
signal result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2337_c7_7acd]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2337_c7_7acd]
signal n8_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2337_c7_7acd]
signal t16_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l2338_c3_1efe]
signal BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2340_c11_c385]
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2340_c7_6b5a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2340_c7_6b5a]
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2340_c7_6b5a]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2340_c7_6b5a]
signal result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2340_c7_6b5a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2340_c7_6b5a]
signal n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2342_c30_f8d0]
signal sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_9f32( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : signed;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.u16_value := ref_toks_7;
      base.sp_relative_shift := ref_toks_8;
      base.is_stack_index_flipped := ref_toks_9;
      base.is_pc_updated := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3
BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_left,
BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_right,
BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d
result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d
result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d
result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d
result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d
result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d
result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d
result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- n8_MUX_uxn_opcodes_h_l2316_c2_753d
n8_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
n8_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
n8_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
n8_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- t16_MUX_uxn_opcodes_h_l2316_c2_753d
t16_MUX_uxn_opcodes_h_l2316_c2_753d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2316_c2_753d_cond,
t16_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue,
t16_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse,
t16_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab
BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_left,
BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_right,
BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75
result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75
result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond,
result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75
result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75
result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond,
result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75
result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output);

-- n8_MUX_uxn_opcodes_h_l2329_c7_cc75
n8_MUX_uxn_opcodes_h_l2329_c7_cc75 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2329_c7_cc75_cond,
n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue,
n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse,
n8_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output);

-- t16_MUX_uxn_opcodes_h_l2329_c7_cc75
t16_MUX_uxn_opcodes_h_l2329_c7_cc75 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2329_c7_cc75_cond,
t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue,
t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse,
t16_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed
BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_left,
BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_right,
BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18
result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18
result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond,
result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18
result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18
result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond,
result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18
result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output);

-- n8_MUX_uxn_opcodes_h_l2332_c7_2c18
n8_MUX_uxn_opcodes_h_l2332_c7_2c18 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2332_c7_2c18_cond,
n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue,
n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse,
n8_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output);

-- t16_MUX_uxn_opcodes_h_l2332_c7_2c18
t16_MUX_uxn_opcodes_h_l2332_c7_2c18 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2332_c7_2c18_cond,
t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue,
t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse,
t16_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output);

-- CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc
CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_x,
CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a
BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_left,
BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_right,
BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd
result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd
result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond,
result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd
result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd
result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond,
result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd
result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output);

-- n8_MUX_uxn_opcodes_h_l2337_c7_7acd
n8_MUX_uxn_opcodes_h_l2337_c7_7acd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2337_c7_7acd_cond,
n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue,
n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse,
n8_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output);

-- t16_MUX_uxn_opcodes_h_l2337_c7_7acd
t16_MUX_uxn_opcodes_h_l2337_c7_7acd : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2337_c7_7acd_cond,
t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue,
t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse,
t16_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe
BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_left,
BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_right,
BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_left,
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_right,
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a
result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a
result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond,
result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output);

-- n8_MUX_uxn_opcodes_h_l2340_c7_6b5a
n8_MUX_uxn_opcodes_h_l2340_c7_6b5a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond,
n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue,
n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse,
n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0
sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_ins,
sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_x,
sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_y,
sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 n8_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 t16_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output,
 n8_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output,
 t16_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output,
 n8_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output,
 t16_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output,
 CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output,
 n8_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output,
 t16_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output,
 BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output,
 n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output,
 sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2326_c3_3828 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2321_c3_2556 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2330_c3_847d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2335_c3_fc1b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2332_c7_2c18_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e3c5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e114_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_99cd_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_a6c8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_2463_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2333_l2338_DUPLICATE_f26f_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9f32_uxn_opcodes_h_l2349_l2311_DUPLICATE_5331_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_right := to_unsigned(3, 2);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2330_c3_847d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2330_c3_847d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_right := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2326_c3_3828 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2326_c3_3828;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2321_c3_2556 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2321_c3_2556;
     VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_y := resize(to_signed(-3, 3), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2335_c3_fc1b := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2335_c3_fc1b;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_left := VAR_phase;
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_left := t16;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse := t16;
     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e114 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e114_return_output := result.u16_value;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2316_c2_753d_return_output := result.is_stack_index_flipped;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2316_c2_753d_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2337_c11_7b3a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2316_c2_753d_return_output := result.is_vram_write;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2333_l2338_DUPLICATE_f26f LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2333_l2338_DUPLICATE_f26f_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2332_c7_2c18_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2316_c6_e0c3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_left;
     BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output := BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e3c5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e3c5_return_output := result.u8_value;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_2463 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_2463_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2340_c11_c385] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_left;
     BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output := BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_a6c8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_a6c8_return_output := result.is_ram_write;

     -- sp_relative_shift[uxn_opcodes_h_l2342_c30_f8d0] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_ins;
     sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_x;
     sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_return_output := sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2329_c11_75ab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_left;
     BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output := BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2332_c11_93ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_99cd LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_99cd_return_output := result.is_opc_done;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2316_c2_753d_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2316_c6_e0c3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2329_c11_75ab_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2332_c11_93ed_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2337_c11_7b3a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_c385_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2333_l2338_DUPLICATE_f26f_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l2333_l2338_DUPLICATE_f26f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_2463_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_2463_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_2463_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_2463_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e114_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e114_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e114_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e114_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e114_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_99cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_99cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_99cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_99cd_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_a6c8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_a6c8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_a6c8_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2332_l2337_l2329_l2340_DUPLICATE_a6c8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e3c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e3c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e3c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e3c5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2316_l2340_l2337_l2332_l2329_DUPLICATE_e3c5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2316_c2_753d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2316_c2_753d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2316_c2_753d_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2316_c2_753d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2332_c7_2c18_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2342_c30_f8d0_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l2334_c3_73cc] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_x <= VAR_CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_return_output := CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l2338_c3_1efe] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_left;
     BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_return_output := BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2340_c7_6b5a] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output := result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2340_c7_6b5a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2340_c7_6b5a] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2340_c7_6b5a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output := result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2340_c7_6b5a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond;
     n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue;
     n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output := n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2340_c7_6b5a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;

     -- Submodule level 2
     VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l2338_c3_1efe_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l2334_c3_73cc_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_6b5a_return_output;
     -- n8_MUX[uxn_opcodes_h_l2337_c7_7acd] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2337_c7_7acd_cond <= VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_cond;
     n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue;
     n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output := n8_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2337_c7_7acd] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output := result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2337_c7_7acd] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;

     -- t16_MUX[uxn_opcodes_h_l2337_c7_7acd] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2337_c7_7acd_cond <= VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_cond;
     t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue;
     t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output := t16_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2337_c7_7acd] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output := result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2337_c7_7acd] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2337_c7_7acd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2329_c7_cc75] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2337_c7_7acd_return_output;
     -- n8_MUX[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2332_c7_2c18_cond <= VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_cond;
     n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue;
     n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output := n8_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;

     -- t16_MUX[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2332_c7_2c18_cond <= VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_cond;
     t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue;
     t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output := t16_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output := result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2332_c7_2c18] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output := result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2332_c7_2c18_return_output;
     -- n8_MUX[uxn_opcodes_h_l2329_c7_cc75] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2329_c7_cc75_cond <= VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_cond;
     n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue;
     n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output := n8_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2329_c7_cc75] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2329_c7_cc75] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output := result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2329_c7_cc75] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2329_c7_cc75] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2329_c7_cc75] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output := result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;

     -- t16_MUX[uxn_opcodes_h_l2329_c7_cc75] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2329_c7_cc75_cond <= VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_cond;
     t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iftrue;
     t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output := t16_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2329_c7_cc75_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     n8_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     n8_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := n8_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- t16_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     t16_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     t16_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := t16_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2316_c2_753d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2316_c2_753d_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_9f32_uxn_opcodes_h_l2349_l2311_DUPLICATE_5331 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9f32_uxn_opcodes_h_l2349_l2311_DUPLICATE_5331_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_9f32(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2316_c2_753d_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2316_c2_753d_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9f32_uxn_opcodes_h_l2349_l2311_DUPLICATE_5331_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_9f32_uxn_opcodes_h_l2349_l2311_DUPLICATE_5331_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
