-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 29
entity sth_0CLK_a9f1e08f is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sth_0CLK_a9f1e08f;
architecture arch of sth_0CLK_a9f1e08f is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2403_c6_eeb5]
signal BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal t8_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2403_c2_4bac]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2416_c11_6884]
signal BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2416_c7_286f]
signal t8_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2416_c7_286f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2416_c7_286f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2416_c7_286f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2416_c7_286f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2416_c7_286f]
signal result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2416_c7_286f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2417_c30_e712]
signal sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2419_c11_a0ab]
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2419_c7_5808]
signal t8_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c7_5808]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c7_5808]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c7_5808]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c7_5808]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2419_c7_5808]
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c7_5808]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_188e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_ram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5
BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_left,
BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_right,
BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output);

-- t8_MUX_uxn_opcodes_h_l2403_c2_4bac
t8_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
t8_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac
result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac
result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac
result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac
result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac
result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac
result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac
result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884
BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_left,
BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_right,
BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output);

-- t8_MUX_uxn_opcodes_h_l2416_c7_286f
t8_MUX_uxn_opcodes_h_l2416_c7_286f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2416_c7_286f_cond,
t8_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue,
t8_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse,
t8_MUX_uxn_opcodes_h_l2416_c7_286f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f
result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f
result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f
result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_cond,
result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f
result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2417_c30_e712
sp_relative_shift_uxn_opcodes_h_l2417_c30_e712 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_ins,
sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_x,
sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_y,
sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab
BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_left,
BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_right,
BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output);

-- t8_MUX_uxn_opcodes_h_l2419_c7_5808
t8_MUX_uxn_opcodes_h_l2419_c7_5808 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2419_c7_5808_cond,
t8_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue,
t8_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse,
t8_MUX_uxn_opcodes_h_l2419_c7_5808_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_cond,
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output,
 t8_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output,
 t8_MUX_uxn_opcodes_h_l2416_c7_286f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_return_output,
 sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output,
 t8_MUX_uxn_opcodes_h_l2419_c7_5808_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2408_c3_0686 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2413_c3_d245 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2424_c3_6652 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2422_c3_564f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2419_c7_5808_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2419_l2403_l2416_DUPLICATE_7cec_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_1920_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_7fb1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_ab58_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_dc7d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2429_l2399_DUPLICATE_6f45_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2422_c3_564f := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2422_c3_564f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2413_c3_d245 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2413_c3_d245;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_right := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2408_c3_0686 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2408_c3_0686;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2424_c3_6652 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2424_c3_6652;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse := t8;
     -- result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d[uxn_opcodes_h_l2419_c7_5808] LATENCY=0
     VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2419_c7_5808_return_output := result.sp_relative_shift;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2416_c11_6884] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_left;
     BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output := BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_dc7d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_dc7d_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_1920 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_1920_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_ab58 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_ab58_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_7fb1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_7fb1_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2403_c6_eeb5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2417_c30_e712] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_ins;
     sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_x;
     sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_return_output := sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2419_l2403_l2416_DUPLICATE_7cec LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2419_l2403_l2416_DUPLICATE_7cec_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2419_c11_a0ab] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_left;
     BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output := BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2403_c6_eeb5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2416_c11_6884_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2419_c11_a0ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_dc7d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_dc7d_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_ab58_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_ab58_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_7fb1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_7fb1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_1920_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2419_l2416_DUPLICATE_1920_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2419_l2403_l2416_DUPLICATE_7cec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2419_l2403_l2416_DUPLICATE_7cec_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2419_l2403_l2416_DUPLICATE_7cec_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2403_c2_4bac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse := VAR_result_sp_relative_shift_FALSE_INPUT_MUX_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2419_c7_5808_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2417_c30_e712_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2419_c7_5808] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2419_c7_5808] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_return_output := result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2419_c7_5808] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2419_c7_5808] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2419_c7_5808] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;

     -- t8_MUX[uxn_opcodes_h_l2419_c7_5808] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2419_c7_5808_cond <= VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_cond;
     t8_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue;
     t8_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_return_output := t8_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2419_c7_5808] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2419_c7_5808_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2416_c7_286f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2416_c7_286f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2416_c7_286f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_return_output := result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2416_c7_286f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;

     -- t8_MUX[uxn_opcodes_h_l2416_c7_286f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2416_c7_286f_cond <= VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_cond;
     t8_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue;
     t8_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_return_output := t8_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2416_c7_286f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2416_c7_286f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2416_c7_286f_return_output;
     -- t8_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := t8_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2403_c2_4bac] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;

     -- Submodule level 4
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2429_l2399_DUPLICATE_6f45 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2429_l2399_DUPLICATE_6f45_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_188e(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2403_c2_4bac_return_output);

     -- Submodule level 5
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2429_l2399_DUPLICATE_6f45_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2429_l2399_DUPLICATE_6f45_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
