-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 40
entity inc2_0CLK_180c5210 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end inc2_0CLK_180c5210;
architecture arch of inc2_0CLK_180c5210 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1378_c6_6e30]
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1378_c2_12d2]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1391_c11_177a]
signal BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1391_c7_f23b]
signal t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1391_c7_f23b]
signal t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1391_c7_f23b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1391_c7_f23b]
signal result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1391_c7_f23b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1391_c7_f23b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1391_c7_f23b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1394_c11_f17b]
signal BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l1394_c7_dd7e]
signal t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1394_c7_dd7e]
signal t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1394_c7_dd7e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1394_c7_dd7e]
signal result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1394_c7_dd7e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1394_c7_dd7e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1394_c7_dd7e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1395_c13_e0fd]
signal BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_return_output : unsigned(8 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1396_c30_871a]
signal sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1401_c11_7c68]
signal BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output : unsigned(0 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l1401_c7_fc9b]
signal t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1401_c7_fc9b]
signal result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1401_c7_fc9b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1401_c7_fc9b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1401_c7_fc9b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1402_c37_0c04]
signal BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1402_c37_e78a]
signal MUX_uxn_opcodes_h_l1402_c37_e78a_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1402_c37_e78a_iftrue : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1402_c37_e78a_iffalse : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1402_c37_e78a_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[uxn_opcodes_h_l1402_c14_e46a]
signal BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_left : unsigned(7 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_return_output : unsigned(8 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_84a2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_vram_write := ref_toks_6;
      base.u8_value := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30
BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_left,
BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_right,
BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2
t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2
t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2
result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2
result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2
result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2
result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a
BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_left,
BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_right,
BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b
t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_cond,
t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue,
t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse,
t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b
t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_cond,
t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue,
t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse,
t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b
result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b
result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b
result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b
BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_left,
BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_right,
BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output);

-- t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e
t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond,
t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue,
t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse,
t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e
t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond,
t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue,
t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse,
t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e
result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e
result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e
result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd
BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_left,
BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_right,
BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1396_c30_871a
sp_relative_shift_uxn_opcodes_h_l1396_c30_871a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_ins,
sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_x,
sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_y,
sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68
BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_left,
BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_right,
BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output);

-- t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b
t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond,
t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue,
t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse,
t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b
result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b
result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04
BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_left,
BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_right,
BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_return_output);

-- MUX_uxn_opcodes_h_l1402_c37_e78a
MUX_uxn_opcodes_h_l1402_c37_e78a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1402_c37_e78a_cond,
MUX_uxn_opcodes_h_l1402_c37_e78a_iftrue,
MUX_uxn_opcodes_h_l1402_c37_e78a_iffalse,
MUX_uxn_opcodes_h_l1402_c37_e78a_return_output);

-- BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a
BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a : entity work.BIN_OP_PLUS_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_left,
BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_right,
BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output,
 t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output,
 t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output,
 t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output,
 t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output,
 t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_return_output,
 sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output,
 t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_return_output,
 MUX_uxn_opcodes_h_l1402_c37_e78a_return_output,
 BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1383_c3_76d3 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1388_c3_a457 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1392_c3_6c24 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_uxn_opcodes_h_l1395_c3_cb3b : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1398_c3_3ecc : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_return_output : unsigned(8 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_uxn_opcodes_h_l1402_c3_de67 : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1403_c3_e26f : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1404_c3_cad2 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1401_c7_fc9b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_left : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_iftrue : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_iffalse : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_return_output : unsigned(8 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1391_l1378_l1401_DUPLICATE_8ebe_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1391_l1394_l1401_DUPLICATE_fbad_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1391_l1401_DUPLICATE_5ce7_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1391_l1394_DUPLICATE_b2e9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1374_l1409_DUPLICATE_071e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1383_c3_76d3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1383_c3_76d3;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1398_c3_3ecc := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1398_c3_3ecc;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_right := to_unsigned(2, 2);
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1404_c3_cad2 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1404_c3_cad2;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_right := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_right := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1403_c3_e26f := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1403_c3_e26f;
     VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1392_c3_6c24 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1392_c3_6c24;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_iffalse := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1388_c3_a457 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1388_c3_a457;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_left := VAR_phase;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_left := VAR_previous_stack_read;
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_left := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse := t16_high;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_left := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse := t16_low;
     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1401_c7_fc9b] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1401_c7_fc9b_return_output := result.stack_address_sp_offset;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l1394_c11_f17b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1391_l1394_DUPLICATE_b2e9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1391_l1394_DUPLICATE_b2e9_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1391_l1378_l1401_DUPLICATE_8ebe LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1391_l1378_l1401_DUPLICATE_8ebe_return_output := result.u8_value;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output := result.is_vram_write;

     -- sp_relative_shift[uxn_opcodes_h_l1396_c30_871a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_ins;
     sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_x;
     sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_return_output := sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1401_c11_7c68] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_left;
     BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output := BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1391_l1401_DUPLICATE_5ce7 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1391_l1401_DUPLICATE_5ce7_return_output := result.sp_relative_shift;

     -- BIN_OP_PLUS[uxn_opcodes_h_l1395_c13_e0fd] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1378_c6_6e30] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_left;
     BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output := BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1391_l1394_l1401_DUPLICATE_fbad LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1391_l1394_l1401_DUPLICATE_fbad_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1391_c11_177a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1402_c37_0c04] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_left;
     BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_return_output := BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1378_c6_6e30_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1391_c11_177a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1394_c11_f17b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1401_c11_7c68_return_output;
     VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1402_c37_0c04_return_output;
     VAR_t16_low_uxn_opcodes_h_l1395_c3_cb3b := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1395_c13_e0fd_return_output, 8);
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1391_l1401_DUPLICATE_5ce7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1391_l1401_DUPLICATE_5ce7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1391_l1394_l1401_DUPLICATE_fbad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1391_l1394_l1401_DUPLICATE_fbad_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1391_l1394_l1401_DUPLICATE_fbad_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1391_l1394_DUPLICATE_b2e9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1391_l1394_DUPLICATE_b2e9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1391_l1378_l1401_DUPLICATE_8ebe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1391_l1378_l1401_DUPLICATE_8ebe_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1391_l1378_l1401_DUPLICATE_8ebe_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1378_c2_12d2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1401_c7_fc9b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1396_c30_871a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue := VAR_t16_low_uxn_opcodes_h_l1395_c3_cb3b;
     VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue := VAR_t16_low_uxn_opcodes_h_l1395_c3_cb3b;
     -- result_is_ram_write_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1401_c7_fc9b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1394_c7_dd7e] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond;
     t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output := t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1401_c7_fc9b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1394_c7_dd7e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;

     -- MUX[uxn_opcodes_h_l1402_c37_e78a] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1402_c37_e78a_cond <= VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_cond;
     MUX_uxn_opcodes_h_l1402_c37_e78a_iftrue <= VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_iftrue;
     MUX_uxn_opcodes_h_l1402_c37_e78a_iffalse <= VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_return_output := MUX_uxn_opcodes_h_l1402_c37_e78a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1401_c7_fc9b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;

     -- Submodule level 2
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_right := VAR_MUX_uxn_opcodes_h_l1402_c37_e78a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;
     -- BIN_OP_PLUS[uxn_opcodes_h_l1402_c14_e46a] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_left <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_left;
     BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_right <= VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_right;
     -- Outputs
     VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_return_output := BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1394_c7_dd7e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1394_c7_dd7e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1391_c7_f23b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1391_c7_f23b] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_cond;
     t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output := t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1394_c7_dd7e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;

     -- Submodule level 3
     VAR_t16_high_uxn_opcodes_h_l1402_c3_de67 := resize(VAR_BIN_OP_PLUS_uxn_opcodes_h_l1402_c14_e46a_return_output, 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue := VAR_t16_high_uxn_opcodes_h_l1402_c3_de67;
     VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue := VAR_t16_high_uxn_opcodes_h_l1402_c3_de67;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1391_c7_f23b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1401_c7_fc9b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1401_c7_fc9b] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_cond;
     t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output := t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1391_c7_f23b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1391_c7_f23b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1401_c7_fc9b_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1394_c7_dd7e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1394_c7_dd7e] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_cond;
     t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output := t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- Submodule level 5
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1394_c7_dd7e_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1391_c7_f23b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1391_c7_f23b] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_cond;
     t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output := t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l1391_c7_f23b_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l1378_c2_12d2] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_cond;
     t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iftrue;
     t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output := t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;

     -- Submodule level 7
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1374_l1409_DUPLICATE_071e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1374_l1409_DUPLICATE_071e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_84a2(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1378_c2_12d2_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1374_l1409_DUPLICATE_071e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_84a2_uxn_opcodes_h_l1374_l1409_DUPLICATE_071e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
