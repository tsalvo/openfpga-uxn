-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity ldz_0CLK_b128164d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_b128164d;
architecture arch of ldz_0CLK_b128164d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_31c4]
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(15 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1437_c2_ef90]
signal t8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_0475]
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1450_c7_ee21]
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_ee21]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1450_c7_ee21]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1450_c7_ee21]
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_ee21]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_ee21]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1450_c7_ee21]
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1450_c7_ee21]
signal t8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1453_c11_1400]
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1453_c7_2903]
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1453_c7_2903]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1453_c7_2903]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : signed(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l1453_c7_2903]
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1453_c7_2903]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1453_c7_2903]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1453_c7_2903]
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1453_c7_2903]
signal t8_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1455_c30_639d]
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1458_c11_3474]
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1458_c7_59ac]
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1458_c7_59ac]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1458_c7_59ac]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1458_c7_59ac]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1458_c7_59ac]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1458_c7_59ac]
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1461_c11_b26b]
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1461_c7_6cf9]
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1461_c7_6cf9]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1461_c7_6cf9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1461_c7_6cf9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1461_c7_6cf9]
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(7 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_e482( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_index_flipped := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.u16_value := ref_toks_4;
      base.is_vram_write := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.is_opc_done := ref_toks_8;
      base.is_ram_write := ref_toks_9;
      base.is_stack_write := ref_toks_10;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_left,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_right,
BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90
tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- t8_MUX_uxn_opcodes_h_l1437_c2_ef90
t8_MUX_uxn_opcodes_h_l1437_c2_ef90 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond,
t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue,
t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse,
t8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_left,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_right,
BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21
tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond,
tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue,
tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse,
tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output);

-- t8_MUX_uxn_opcodes_h_l1450_c7_ee21
t8_MUX_uxn_opcodes_h_l1450_c7_ee21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond,
t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue,
t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse,
t8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_left,
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_right,
BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1453_c7_2903
tmp8_MUX_uxn_opcodes_h_l1453_c7_2903 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_cond,
tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue,
tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse,
tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output);

-- t8_MUX_uxn_opcodes_h_l1453_c7_2903
t8_MUX_uxn_opcodes_h_l1453_c7_2903 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1453_c7_2903_cond,
t8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue,
t8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse,
t8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1455_c30_639d
sp_relative_shift_uxn_opcodes_h_l1455_c30_639d : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_ins,
sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_x,
sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_y,
sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_left,
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_right,
BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_cond,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac
tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_cond,
tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue,
tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse,
tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_left,
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_right,
BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9
tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond,
tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue,
tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse,
tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 t8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output,
 tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output,
 t8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_return_output,
 tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output,
 t8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output,
 sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output,
 tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output,
 tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_1392 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_2f77 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_94cf : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_return_output : signed(3 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_c57b_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_aa0c : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_da4e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1437_l1461_l1458_l1453_l1450_DUPLICATE_9ef4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_d00d_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_2e8f_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_c709_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_9c54_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_2472_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1469_l1433_DUPLICATE_8a99_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_x := signed(std_logic_vector(resize(to_unsigned(1, 1), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_1392 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1447_c3_1392;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_94cf := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1451_c3_94cf;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_da4e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1464_c3_da4e;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_aa0c := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1459_c3_aa0c;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_right := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_2f77 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1442_c3_2f77;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_left := VAR_phase;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse := tmp8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1437_l1461_l1458_l1453_l1450_DUPLICATE_9ef4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1437_l1461_l1458_l1453_l1450_DUPLICATE_9ef4_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1437_c6_31c4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_left;
     BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output := BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_9c54 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_9c54_return_output := result.is_stack_write;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1456_c22_c57b] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_c57b_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_c709 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_c709_return_output := result.is_opc_done;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1450_c11_0475] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_left;
     BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output := BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1458_c11_3474] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_left;
     BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output := BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_2472 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_2472_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l1455_c30_639d] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_ins;
     sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_x;
     sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_return_output := sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l1453_c11_1400] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_left;
     BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output := BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1461_c11_b26b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_2e8f LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_2e8f_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_d00d LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_d00d_return_output := result.u16_value;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1437_c6_31c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1450_c11_0475_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1453_c11_1400_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1458_c11_3474_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1461_c11_b26b_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1456_c22_c57b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_2e8f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1458_l1450_DUPLICATE_2e8f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_d00d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_d00d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l1437_l1450_l1453_DUPLICATE_d00d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_c709_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_c709_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_c709_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_c709_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_9c54_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_9c54_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_9c54_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1458_l1450_l1461_l1453_DUPLICATE_9c54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_2472_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_2472_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1458_l1461_l1453_DUPLICATE_2472_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1437_l1461_l1458_l1453_l1450_DUPLICATE_9ef4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1437_l1461_l1458_l1453_l1450_DUPLICATE_9ef4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1437_l1461_l1458_l1453_l1450_DUPLICATE_9ef4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1437_l1461_l1458_l1453_l1450_DUPLICATE_9ef4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1437_l1461_l1458_l1453_l1450_DUPLICATE_9ef4_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1437_c2_ef90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1455_c30_639d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1461_c7_6cf9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1461_c7_6cf9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1458_c7_59ac] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1461_c7_6cf9] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1453_c7_2903] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output := result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1461_c7_6cf9] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond;
     tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output := tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;

     -- t8_MUX[uxn_opcodes_h_l1453_c7_2903] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1453_c7_2903_cond <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_cond;
     t8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue;
     t8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output := t8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1461_c7_6cf9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output := result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1461_c7_6cf9_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1458_c7_59ac] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;

     -- t8_MUX[uxn_opcodes_h_l1450_c7_ee21] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond;
     t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue;
     t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output := t8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1458_c7_59ac] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output := result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1458_c7_59ac] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_cond;
     tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output := tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1453_c7_2903] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1450_c7_ee21] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output := result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1458_c7_59ac] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1458_c7_59ac] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1458_c7_59ac_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1450_c7_ee21] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1453_c7_2903] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output := result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1453_c7_2903] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1453_c7_2903] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1453_c7_2903] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1453_c7_2903] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_cond;
     tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output := tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;

     -- t8_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := t8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1453_c7_2903_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1450_c7_ee21] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output := result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1450_c7_ee21] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1450_c7_ee21] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1450_c7_ee21] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_cond;
     tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output := tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1450_c7_ee21] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1450_c7_ee21_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1437_c2_ef90] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;

     -- Submodule level 6
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1469_l1433_DUPLICATE_8a99 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1469_l1433_DUPLICATE_8a99_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e482(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1437_c2_ef90_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1469_l1433_DUPLICATE_8a99_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e482_uxn_opcodes_h_l1469_l1433_DUPLICATE_8a99_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
