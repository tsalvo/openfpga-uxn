-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity sub_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_bacf6a1d;
architecture arch of sub_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2335_c6_247d]
signal BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2335_c1_35bd]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2335_c2_6d8d]
signal n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2335_c2_6d8d]
signal t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2335_c2_6d8d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2335_c2_6d8d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2335_c2_6d8d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2335_c2_6d8d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2335_c2_6d8d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2335_c2_6d8d]
signal result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l2336_c3_f0d1[uxn_opcodes_h_l2336_c3_f0d1]
signal printf_uxn_opcodes_h_l2336_c3_f0d1_uxn_opcodes_h_l2336_c3_f0d1_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2340_c11_eb48]
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2340_c7_cceb]
signal n8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2340_c7_cceb]
signal t8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2340_c7_cceb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2340_c7_cceb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2340_c7_cceb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2340_c7_cceb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2340_c7_cceb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2340_c7_cceb]
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2343_c11_db2b]
signal BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2343_c7_3d8e]
signal n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2343_c7_3d8e]
signal t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2343_c7_3d8e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2343_c7_3d8e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2343_c7_3d8e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2343_c7_3d8e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2343_c7_3d8e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2343_c7_3d8e]
signal result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2346_c11_4a71]
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2346_c7_e36c]
signal n8_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2346_c7_e36c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2346_c7_e36c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2346_c7_e36c]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2346_c7_e36c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2346_c7_e36c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2346_c7_e36c]
signal result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2349_c30_8610]
signal sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2352_c21_9278]
signal BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2354_c11_e8d6]
signal BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2354_c7_b62e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2354_c7_b62e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2354_c7_b62e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4e73( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d
BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_left,
BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_right,
BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_return_output);

-- n8_MUX_uxn_opcodes_h_l2335_c2_6d8d
n8_MUX_uxn_opcodes_h_l2335_c2_6d8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond,
n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue,
n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse,
n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

-- t8_MUX_uxn_opcodes_h_l2335_c2_6d8d
t8_MUX_uxn_opcodes_h_l2335_c2_6d8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond,
t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue,
t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse,
t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

-- printf_uxn_opcodes_h_l2336_c3_f0d1_uxn_opcodes_h_l2336_c3_f0d1
printf_uxn_opcodes_h_l2336_c3_f0d1_uxn_opcodes_h_l2336_c3_f0d1 : entity work.printf_uxn_opcodes_h_l2336_c3_f0d1_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l2336_c3_f0d1_uxn_opcodes_h_l2336_c3_f0d1_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_left,
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_right,
BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output);

-- n8_MUX_uxn_opcodes_h_l2340_c7_cceb
n8_MUX_uxn_opcodes_h_l2340_c7_cceb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond,
n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue,
n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse,
n8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output);

-- t8_MUX_uxn_opcodes_h_l2340_c7_cceb
t8_MUX_uxn_opcodes_h_l2340_c7_cceb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond,
t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue,
t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse,
t8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_cond,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b
BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_left,
BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_right,
BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output);

-- n8_MUX_uxn_opcodes_h_l2343_c7_3d8e
n8_MUX_uxn_opcodes_h_l2343_c7_3d8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond,
n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue,
n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse,
n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output);

-- t8_MUX_uxn_opcodes_h_l2343_c7_3d8e
t8_MUX_uxn_opcodes_h_l2343_c7_3d8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond,
t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue,
t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse,
t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_left,
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_right,
BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output);

-- n8_MUX_uxn_opcodes_h_l2346_c7_e36c
n8_MUX_uxn_opcodes_h_l2346_c7_e36c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2346_c7_e36c_cond,
n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue,
n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse,
n8_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2349_c30_8610
sp_relative_shift_uxn_opcodes_h_l2349_c30_8610 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_ins,
sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_x,
sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_y,
sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278
BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_left,
BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_right,
BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6
BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_left,
BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_right,
BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_return_output,
 n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
 t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output,
 n8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output,
 t8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output,
 n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output,
 t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output,
 n8_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output,
 sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2337_c3_7279 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l2336_c3_f0d1_uxn_opcodes_h_l2336_c3_f0d1_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2341_c3_cf09 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2351_c3_3d3f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_252b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_86c4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_c200_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_6319_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2346_l2340_l2354_l2343_DUPLICATE_2145_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2346_l2343_DUPLICATE_7640_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2360_l2331_DUPLICATE_9bdd_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2341_c3_cf09 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2341_c3_cf09;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2337_c3_7279 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2337_c3_7279;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2351_c3_3d3f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2351_c3_3d3f;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_right := to_unsigned(2, 2);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2346_l2340_l2354_l2343_DUPLICATE_2145 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2346_l2340_l2354_l2343_DUPLICATE_2145_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2335_c6_247d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_left;
     BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output := BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2343_c11_db2b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_left;
     BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output := BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2340_c11_eb48] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_left;
     BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output := BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2346_l2343_DUPLICATE_7640 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2346_l2343_DUPLICATE_7640_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2346_c11_4a71] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_left;
     BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output := BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2349_c30_8610] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_ins;
     sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_x;
     sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_return_output := sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_return_output;

     -- BIN_OP_MINUS[uxn_opcodes_h_l2352_c21_9278] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_c200 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_c200_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2354_c11_e8d6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_252b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_252b_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_6319 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_6319_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_86c4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_86c4_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2335_c6_247d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2340_c11_eb48_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2343_c11_db2b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2346_c11_4a71_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2354_c11_e8d6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2352_c21_9278_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_c200_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_c200_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_c200_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_c200_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2346_l2340_l2354_l2343_DUPLICATE_2145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2346_l2340_l2354_l2343_DUPLICATE_2145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2346_l2340_l2354_l2343_DUPLICATE_2145_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2346_l2340_l2354_l2343_DUPLICATE_2145_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_86c4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_86c4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_86c4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_86c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_252b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_252b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_252b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2335_l2340_l2354_l2343_DUPLICATE_252b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2346_l2343_DUPLICATE_7640_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2346_l2343_DUPLICATE_7640_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_6319_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_6319_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_6319_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2335_l2346_l2340_l2343_DUPLICATE_6319_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2349_c30_8610_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2354_c7_b62e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output;

     -- t8_MUX[uxn_opcodes_h_l2343_c7_3d8e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond <= VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond;
     t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue;
     t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output := t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l2335_c1_35bd] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2354_c7_b62e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2354_c7_b62e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2346_c7_e36c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2346_c7_e36c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_cond;
     n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue;
     n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output := n8_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2346_c7_e36c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2346_c7_e36c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2346_c7_e36c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l2336_c3_f0d1_uxn_opcodes_h_l2336_c3_f0d1_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l2335_c1_35bd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2354_c7_b62e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2346_c7_e36c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2343_c7_3d8e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2346_c7_e36c] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2343_c7_3d8e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2346_c7_e36c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;

     -- t8_MUX[uxn_opcodes_h_l2340_c7_cceb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond <= VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond;
     t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue;
     t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output := t8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;

     -- n8_MUX[uxn_opcodes_h_l2343_c7_3d8e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond <= VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond;
     n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue;
     n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output := n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2343_c7_3d8e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;

     -- printf_uxn_opcodes_h_l2336_c3_f0d1[uxn_opcodes_h_l2336_c3_f0d1] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l2336_c3_f0d1_uxn_opcodes_h_l2336_c3_f0d1_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l2336_c3_f0d1_uxn_opcodes_h_l2336_c3_f0d1_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2346_c7_e36c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2340_c7_cceb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2343_c7_3d8e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;

     -- t8_MUX[uxn_opcodes_h_l2335_c2_6d8d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond <= VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond;
     t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue;
     t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output := t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2340_c7_cceb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2343_c7_3d8e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;

     -- n8_MUX[uxn_opcodes_h_l2340_c7_cceb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_cond;
     n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue;
     n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output := n8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2340_c7_cceb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output := result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2343_c7_3d8e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2343_c7_3d8e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2340_c7_cceb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2335_c2_6d8d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2340_c7_cceb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2335_c2_6d8d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2340_c7_cceb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;

     -- n8_MUX[uxn_opcodes_h_l2335_c2_6d8d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond;
     n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue;
     n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output := n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2335_c2_6d8d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2340_c7_cceb_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2335_c2_6d8d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2335_c2_6d8d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2335_c2_6d8d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2360_l2331_DUPLICATE_9bdd LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2360_l2331_DUPLICATE_9bdd_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4e73(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2335_c2_6d8d_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2360_l2331_DUPLICATE_9bdd_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4e73_uxn_opcodes_h_l2360_l2331_DUPLICATE_9bdd_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
