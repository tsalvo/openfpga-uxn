-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity sta_0CLK_9159c4aa is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end sta_0CLK_9159c4aa;
architecture arch of sta_0CLK_9159c4aa is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2070_c6_e731]
signal BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal n8_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2070_c2_6e26]
signal t16_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2078_c11_c43f]
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal n8_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2078_c7_7c67]
signal t16_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2082_c11_8650]
signal BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2082_c7_dae9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2082_c7_dae9]
signal result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2082_c7_dae9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2082_c7_dae9]
signal result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2082_c7_dae9]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : signed(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2082_c7_dae9]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2082_c7_dae9]
signal n8_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(7 downto 0);

-- t16_MUX[uxn_opcodes_h_l2082_c7_dae9]
signal t16_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2085_c30_4efa]
signal sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2087_c11_4012]
signal BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2087_c7_5385]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2087_c7_5385]
signal result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2087_c7_5385]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2087_c7_5385]
signal result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2087_c7_5385]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2087_c7_5385]
signal n8_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2094_c11_0524]
signal BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2094_c7_f178]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2094_c7_f178]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_return_output : unsigned(0 downto 0);

function CAST_TO_uint8_t_uint16_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(15 downto 0);
  variable return_output : unsigned(7 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,8)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.u8_value := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.is_stack_operation_16bit := ref_toks_7;
      base.is_ram_write := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731
BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_left,
BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_right,
BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26
result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26
result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26
result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26
result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26
result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26
result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- n8_MUX_uxn_opcodes_h_l2070_c2_6e26
n8_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
n8_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- t16_MUX_uxn_opcodes_h_l2070_c2_6e26
t16_MUX_uxn_opcodes_h_l2070_c2_6e26 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2070_c2_6e26_cond,
t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue,
t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse,
t16_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f
BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_left,
BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_right,
BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67
result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67
result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67
result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- n8_MUX_uxn_opcodes_h_l2078_c7_7c67
n8_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
n8_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- t16_MUX_uxn_opcodes_h_l2078_c7_7c67
t16_MUX_uxn_opcodes_h_l2078_c7_7c67 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2078_c7_7c67_cond,
t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue,
t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse,
t16_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650
BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_left,
BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_right,
BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9
result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9
result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond,
result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9
result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9
result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond,
result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9
result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9
result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output);

-- n8_MUX_uxn_opcodes_h_l2082_c7_dae9
n8_MUX_uxn_opcodes_h_l2082_c7_dae9 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2082_c7_dae9_cond,
n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue,
n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse,
n8_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output);

-- t16_MUX_uxn_opcodes_h_l2082_c7_dae9
t16_MUX_uxn_opcodes_h_l2082_c7_dae9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2082_c7_dae9_cond,
t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue,
t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse,
t16_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa
sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_ins,
sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_x,
sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_y,
sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012
BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_left,
BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_right,
BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385
result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385
result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond,
result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385
result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385
result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond,
result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385
result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_return_output);

-- n8_MUX_uxn_opcodes_h_l2087_c7_5385
n8_MUX_uxn_opcodes_h_l2087_c7_5385 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2087_c7_5385_cond,
n8_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue,
n8_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse,
n8_MUX_uxn_opcodes_h_l2087_c7_5385_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524
BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_left,
BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_right,
BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178
result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 n8_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 t16_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 n8_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 t16_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output,
 n8_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output,
 t16_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output,
 sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_return_output,
 n8_MUX_uxn_opcodes_h_l2087_c7_5385_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2075_c3_31ec : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2080_c3_9d0d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2078_c7_7c67_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2088_c8_eb99_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_cc83_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_1fbc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2082_l2070_l2078_DUPLICATE_5abd_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2070_l2087_l2078_DUPLICATE_8ba2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2082_l2070_l2078_l2094_DUPLICATE_63ee_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2082_l2087_l2078_l2094_DUPLICATE_fb89_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2099_l2065_DUPLICATE_fe52_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_y := resize(to_signed(-3, 3), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2075_c3_31ec := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2075_c3_31ec;
     VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_right := to_unsigned(4, 3);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2080_c3_9d0d := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2080_c3_9d0d;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_left := VAR_phase;
     VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2082_l2087_l2078_l2094_DUPLICATE_fb89 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2082_l2087_l2078_l2094_DUPLICATE_fb89_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2094_c11_0524] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_left;
     BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_return_output := BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2078_c7_7c67_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2087_c11_4012] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_left;
     BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output := BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2085_c30_4efa] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_ins;
     sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_x;
     sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_return_output := sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_1fbc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_1fbc_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2082_c11_8650] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_left;
     BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output := BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_cc83 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_cc83_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2070_c6_e731] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_left;
     BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output := BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;

     -- CAST_TO_uint8_t[uxn_opcodes_h_l2088_c8_eb99] LATENCY=0
     VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2088_c8_eb99_return_output := CAST_TO_uint8_t_uint16_t(
     VAR_previous_stack_read);

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2070_l2087_l2078_DUPLICATE_8ba2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2070_l2087_l2078_DUPLICATE_8ba2_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2082_l2070_l2078_DUPLICATE_5abd LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2082_l2070_l2078_DUPLICATE_5abd_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2078_c11_c43f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_left;
     BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output := BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2082_l2070_l2078_l2094_DUPLICATE_63ee LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2082_l2070_l2078_l2094_DUPLICATE_63ee_return_output := result.is_ram_write;

     -- result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2078_c7_7c67_return_output := result.is_stack_operation_16bit;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2070_c6_e731_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2078_c11_c43f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2082_c11_8650_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2087_c11_4012_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2094_c11_0524_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2088_c8_eb99_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue := VAR_CAST_TO_uint8_t_uxn_opcodes_h_l2088_c8_eb99_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2082_l2070_l2078_DUPLICATE_5abd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2082_l2070_l2078_DUPLICATE_5abd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2082_l2070_l2078_DUPLICATE_5abd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_cc83_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_cc83_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_cc83_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_cc83_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2082_l2087_l2078_l2094_DUPLICATE_fb89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2082_l2087_l2078_l2094_DUPLICATE_fb89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2082_l2087_l2078_l2094_DUPLICATE_fb89_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2082_l2087_l2078_l2094_DUPLICATE_fb89_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2082_l2070_l2078_l2094_DUPLICATE_63ee_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2082_l2070_l2078_l2094_DUPLICATE_63ee_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2082_l2070_l2078_l2094_DUPLICATE_63ee_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2082_l2070_l2078_l2094_DUPLICATE_63ee_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2070_l2087_l2078_DUPLICATE_8ba2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2070_l2087_l2078_DUPLICATE_8ba2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2070_l2087_l2078_DUPLICATE_8ba2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_1fbc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_1fbc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_1fbc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2082_l2070_l2087_l2078_DUPLICATE_1fbc_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_result_is_stack_operation_16bit_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2085_c30_4efa_return_output;
     -- n8_MUX[uxn_opcodes_h_l2087_c7_5385] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2087_c7_5385_cond <= VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_cond;
     n8_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue;
     n8_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_return_output := n8_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2094_c7_f178] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_return_output;

     -- t16_MUX[uxn_opcodes_h_l2082_c7_dae9] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2082_c7_dae9_cond <= VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_cond;
     t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue;
     t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output := t16_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2087_c7_5385] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2087_c7_5385] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output := result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2082_c7_dae9] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2094_c7_f178] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2087_c7_5385] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output := result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2094_c7_f178_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2094_c7_f178_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2082_c7_dae9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output := result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;

     -- t16_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := t16_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2087_c7_5385] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2082_c7_dae9] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output := result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2082_c7_dae9] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2082_c7_dae9_cond <= VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_cond;
     n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue;
     n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output := n8_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2087_c7_5385] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2082_c7_dae9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2087_c7_5385_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2082_c7_dae9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;

     -- n8_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := n8_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- t16_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := t16_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2082_c7_dae9] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2082_c7_dae9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;
     -- n8_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := n8_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2078_c7_7c67] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse := VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2078_c7_7c67_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2070_c2_6e26] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2099_l2065_DUPLICATE_fe52 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2099_l2065_DUPLICATE_fe52_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2070_c2_6e26_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2099_l2065_DUPLICATE_fe52_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c7f2_uxn_opcodes_h_l2099_l2065_DUPLICATE_fe52_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
