-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 67
entity swp2_0CLK_814c2afd is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end swp2_0CLK_814c2afd;
architecture arch of swp2_0CLK_814c2afd is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n16_high : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n16_low : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16_high : unsigned(7 downto 0);
signal REG_COMB_t16_low : unsigned(7 downto 0);
signal REG_COMB_n16_high : unsigned(7 downto 0);
signal REG_COMB_n16_low : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2602_c6_90b0]
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2602_c2_dc54]
signal t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2615_c11_ef1e]
signal BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(0 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2615_c7_a7ed]
signal t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2618_c11_a574]
signal BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(0 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);

-- t16_high_MUX[uxn_opcodes_h_l2618_c7_b0cc]
signal t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
signal t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2622_c11_70b1]
signal BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output : unsigned(0 downto 0);

-- t16_low_MUX[uxn_opcodes_h_l2622_c7_7d8c]
signal t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(7 downto 0);
signal t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(7 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2622_c7_7d8c]
signal n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2622_c7_7d8c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2622_c7_7d8c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2622_c7_7d8c]
signal result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2622_c7_7d8c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2622_c7_7d8c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(0 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2622_c7_7d8c]
signal n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2626_c11_48f2]
signal BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output : unsigned(0 downto 0);

-- n16_high_MUX[uxn_opcodes_h_l2626_c7_df69]
signal n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(7 downto 0);
signal n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2626_c7_df69]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2626_c7_df69]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2626_c7_df69]
signal result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2626_c7_df69]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2626_c7_df69]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(0 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2626_c7_df69]
signal n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2628_c30_c091]
signal sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2633_c11_207a]
signal BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2633_c7_7995]
signal result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2633_c7_7995]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2633_c7_7995]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2633_c7_7995]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : unsigned(3 downto 0);

-- n16_low_MUX[uxn_opcodes_h_l2633_c7_7995]
signal n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : unsigned(7 downto 0);
signal n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2639_c11_047e]
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2639_c7_407e]
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c7_407e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c7_407e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_return_output : unsigned(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2643_c11_037c]
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2643_c7_3154]
signal result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2643_c7_3154]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2643_c7_3154]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_return_output : unsigned(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a47b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0
BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_left,
BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_right,
BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54
t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54
n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54
result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54
result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54
result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54
n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54
t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond,
t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue,
t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse,
t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e
BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_left,
BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_right,
BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed
t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed
n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed
result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed
result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed
result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed
result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed
n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed
t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond,
t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue,
t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse,
t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574
BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_left,
BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_right,
BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc
t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc
n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc
result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc
result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc
n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc
t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond,
t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue,
t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse,
t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1
BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_left,
BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_right,
BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output);

-- t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c
t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond,
t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue,
t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse,
t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c
n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond,
n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue,
n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse,
n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c
result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c
n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond,
n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue,
n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse,
n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2
BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_left,
BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_right,
BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output);

-- n16_high_MUX_uxn_opcodes_h_l2626_c7_df69
n16_high_MUX_uxn_opcodes_h_l2626_c7_df69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_cond,
n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue,
n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse,
n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69
result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69
result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69
result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_cond,
result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69
result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2626_c7_df69
n16_low_MUX_uxn_opcodes_h_l2626_c7_df69 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_cond,
n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue,
n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse,
n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2628_c30_c091
sp_relative_shift_uxn_opcodes_h_l2628_c30_c091 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_ins,
sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_x,
sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_y,
sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a
BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_left,
BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_right,
BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995
result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_cond,
result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995
result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995
result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_return_output);

-- n16_low_MUX_uxn_opcodes_h_l2633_c7_7995
n16_low_MUX_uxn_opcodes_h_l2633_c7_7995 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_cond,
n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue,
n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse,
n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e
BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_left,
BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_right,
BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e
result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_cond,
result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_left,
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_right,
BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_cond,
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16_high,
 t16_low,
 n16_high,
 n16_low,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output,
 t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output,
 t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output,
 t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output,
 t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output,
 n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output,
 n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output,
 n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_return_output,
 n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_return_output,
 sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_return_output,
 n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2607_c3_9708 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2612_c3_931b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2616_c3_e69d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2620_c3_8319 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse : unsigned(7 downto 0);
 variable VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output : unsigned(0 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(7 downto 0);
 variable VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2624_c3_5182 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output : unsigned(0 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(7 downto 0);
 variable VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2630_c3_789a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_return_output : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2635_c3_ce46 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2636_c3_14e1 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse : unsigned(7 downto 0);
 variable VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_8f85 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2644_c3_1c35 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2643_c7_3154_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2602_l2622_DUPLICATE_c568_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2618_l2633_l2622_l2615_DUPLICATE_b636_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2626_l2618_l2622_l2615_DUPLICATE_c74f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2598_l2649_DUPLICATE_7654_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16_high : unsigned(7 downto 0);
variable REG_VAR_t16_low : unsigned(7 downto 0);
variable REG_VAR_n16_high : unsigned(7 downto 0);
variable REG_VAR_n16_low : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16_high := t16_high;
  REG_VAR_t16_low := t16_low;
  REG_VAR_n16_high := n16_high;
  REG_VAR_n16_low := n16_low;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2636_c3_14e1 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2636_c3_14e1;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2630_c3_789a := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2630_c3_789a;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2620_c3_8319 := resize(to_unsigned(4, 3), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2620_c3_8319;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_x := signed(std_logic_vector(resize(to_unsigned(4, 3), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_right := to_unsigned(3, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2635_c3_ce46 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2635_c3_ce46;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2616_c3_e69d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2616_c3_e69d;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2607_c3_9708 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2607_c3_9708;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2624_c3_5182 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2624_c3_5182;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := to_unsigned(0, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2612_c3_931b := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2612_c3_931b;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_right := to_unsigned(7, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2644_c3_1c35 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2644_c3_1c35;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_8f85 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2640_c3_8f85;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_right := to_unsigned(6, 3);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_ins := VAR_ins;
     VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue := n16_high;
     VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse := n16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue := n16_high;
     VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue := n16_low;
     VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse := n16_low;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue := n16_low;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_left := VAR_phase;
     VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue := VAR_previous_stack_read;
     VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue := VAR_previous_stack_read;
     VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := VAR_previous_stack_read;
     VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := t16_high;
     VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := t16_high;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := t16_low;
     VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse := t16_low;
     -- sp_relative_shift[uxn_opcodes_h_l2628_c30_c091] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_ins;
     sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_x;
     sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_return_output := sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2618_l2633_l2622_l2615_DUPLICATE_b636 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2618_l2633_l2622_l2615_DUPLICATE_b636_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2602_c6_90b0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_left;
     BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output := BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2615_c11_ef1e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2643_c7_3154] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2643_c7_3154_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2626_l2618_l2622_l2615_DUPLICATE_c74f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2626_l2618_l2622_l2615_DUPLICATE_c74f_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2633_c11_207a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output := result.is_vram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2643_c11_037c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output := result.is_ram_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2602_l2622_DUPLICATE_c568 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2602_l2622_DUPLICATE_c568_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output := result.is_pc_updated;

     -- BIN_OP_EQ[uxn_opcodes_h_l2639_c11_047e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_left;
     BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output := BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2618_c11_a574] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_left;
     BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output := BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2626_c11_48f2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output := result.is_stack_index_flipped;

     -- BIN_OP_EQ[uxn_opcodes_h_l2622_c11_70b1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_left;
     BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output := BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;

     -- Submodule level 1
     VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2602_c6_90b0_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2615_c11_ef1e_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2618_c11_a574_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2622_c11_70b1_return_output;
     VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2626_c11_48f2_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2633_c11_207a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2639_c11_047e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2643_c11_037c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2618_l2633_l2622_l2615_DUPLICATE_b636_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2618_l2633_l2622_l2615_DUPLICATE_b636_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2618_l2633_l2622_l2615_DUPLICATE_b636_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2618_l2633_l2622_l2615_DUPLICATE_b636_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2639_l2633_l2626_l2622_DUPLICATE_dfe8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2626_l2618_l2622_l2615_DUPLICATE_c74f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2626_l2618_l2622_l2615_DUPLICATE_c74f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2626_l2618_l2622_l2615_DUPLICATE_c74f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2626_l2618_l2622_l2615_DUPLICATE_c74f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2602_l2622_DUPLICATE_c568_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2602_l2622_DUPLICATE_c568_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2602_l2622_DUPLICATE_c568_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2602_l2622_DUPLICATE_c568_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2618_l2615_l2643_l2602_l2622_DUPLICATE_c568_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2602_c2_dc54_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2643_c7_3154_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2628_c30_c091_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2643_c7_3154] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2643_c7_3154] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2633_c7_7995] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_cond;
     n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_return_output := n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2633_c7_7995] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2626_c7_df69] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2643_c7_3154] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_return_output := result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l2626_c7_df69] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_cond;
     n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_return_output := n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2622_c7_7d8c] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond;
     t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output := t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- Submodule level 2
     VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2643_c7_3154_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2643_c7_3154_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2643_c7_3154_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2639_c7_407e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l2622_c7_7d8c] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond;
     n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output := n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2622_c7_7d8c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2626_c7_df69] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2626_c7_df69] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_cond;
     n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_return_output := n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2639_c7_407e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_return_output := result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2639_c7_407e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_return_output;

     -- Submodule level 3
     VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2639_c7_407e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2639_c7_407e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2639_c7_407e_return_output;
     VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_t16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     -- n16_high_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2633_c7_7995] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_return_output := result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2622_c7_7d8c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2622_c7_7d8c] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond;
     n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output := n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;

     -- t16_high_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2633_c7_7995] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2633_c7_7995] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;

     -- Submodule level 4
     VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2633_c7_7995_return_output;
     REG_VAR_t16_high := VAR_t16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;
     VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_t16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     -- n16_low_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- t16_low_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2626_c7_df69] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_return_output := result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2626_c7_df69] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2626_c7_df69] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- Submodule level 5
     VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_n16_high_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2626_c7_df69_return_output;
     REG_VAR_t16_low := VAR_t16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;
     -- n16_low_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- n16_high_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2622_c7_7d8c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2622_c7_7d8c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2622_c7_7d8c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;

     -- Submodule level 6
     REG_VAR_n16_high := VAR_n16_high_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;
     VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_n16_low_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2622_c7_7d8c_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2618_c7_b0cc] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;

     -- n16_low_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- Submodule level 7
     REG_VAR_n16_low := VAR_n16_low_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2618_c7_b0cc_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2615_c7_a7ed] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;

     -- Submodule level 8
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2615_c7_a7ed_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2602_c2_dc54] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output;

     -- Submodule level 9
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2598_l2649_DUPLICATE_7654 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2598_l2649_DUPLICATE_7654_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a47b(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2602_c2_dc54_return_output);

     -- Submodule level 10
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2598_l2649_DUPLICATE_7654_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l2598_l2649_DUPLICATE_7654_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16_high <= REG_VAR_t16_high;
REG_COMB_t16_low <= REG_VAR_t16_low;
REG_COMB_n16_high <= REG_VAR_n16_high;
REG_COMB_n16_low <= REG_VAR_n16_low;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16_high <= REG_COMB_t16_high;
     t16_low <= REG_COMB_t16_low;
     n16_high <= REG_COMB_n16_high;
     n16_low <= REG_COMB_n16_low;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
