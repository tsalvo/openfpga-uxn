-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity equ_0CLK_7883ef49 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_7883ef49;
architecture arch of equ_0CLK_7883ef49 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1140_c6_b37c]
signal BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1140_c2_aa8c]
signal n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1140_c2_aa8c]
signal result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1140_c2_aa8c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1140_c2_aa8c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1140_c2_aa8c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1140_c2_aa8c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1140_c2_aa8c]
signal t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1147_c11_c3d5]
signal BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1147_c7_b81b]
signal n8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1147_c7_b81b]
signal result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1147_c7_b81b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1147_c7_b81b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1147_c7_b81b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1147_c7_b81b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1147_c7_b81b]
signal t8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1150_c11_0dd1]
signal BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1150_c7_a553]
signal n8_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1150_c7_a553]
signal result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1150_c7_a553]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1150_c7_a553]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1150_c7_a553]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1150_c7_a553]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1150_c7_a553]
signal t8_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1153_c11_b258]
signal BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1153_c7_76c0]
signal n8_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1153_c7_76c0]
signal result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1153_c7_76c0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1153_c7_76c0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1153_c7_76c0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1153_c7_76c0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1156_c30_890f]
signal sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1159_c21_06c1]
signal BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1159_c21_dcf2]
signal MUX_uxn_opcodes_h_l1159_c21_dcf2_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1159_c21_dcf2_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1159_c21_dcf2_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1159_c21_dcf2_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1161_c11_eade]
signal BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1161_c7_49ca]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1161_c7_49ca]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1161_c7_49ca]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c
BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_left,
BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_right,
BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output);

-- n8_MUX_uxn_opcodes_h_l1140_c2_aa8c
n8_MUX_uxn_opcodes_h_l1140_c2_aa8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond,
n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue,
n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse,
n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c
result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c
result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c
result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output);

-- t8_MUX_uxn_opcodes_h_l1140_c2_aa8c
t8_MUX_uxn_opcodes_h_l1140_c2_aa8c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond,
t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue,
t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse,
t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5
BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_left,
BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_right,
BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output);

-- n8_MUX_uxn_opcodes_h_l1147_c7_b81b
n8_MUX_uxn_opcodes_h_l1147_c7_b81b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond,
n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue,
n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse,
n8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b
result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b
result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b
result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output);

-- t8_MUX_uxn_opcodes_h_l1147_c7_b81b
t8_MUX_uxn_opcodes_h_l1147_c7_b81b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond,
t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue,
t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse,
t8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1
BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_left,
BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_right,
BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output);

-- n8_MUX_uxn_opcodes_h_l1150_c7_a553
n8_MUX_uxn_opcodes_h_l1150_c7_a553 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1150_c7_a553_cond,
n8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue,
n8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse,
n8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_cond,
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_return_output);

-- t8_MUX_uxn_opcodes_h_l1150_c7_a553
t8_MUX_uxn_opcodes_h_l1150_c7_a553 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1150_c7_a553_cond,
t8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue,
t8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse,
t8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258
BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_left,
BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_right,
BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output);

-- n8_MUX_uxn_opcodes_h_l1153_c7_76c0
n8_MUX_uxn_opcodes_h_l1153_c7_76c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1153_c7_76c0_cond,
n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue,
n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse,
n8_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1156_c30_890f
sp_relative_shift_uxn_opcodes_h_l1156_c30_890f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_ins,
sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_x,
sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_y,
sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1
BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_left,
BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_right,
BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_return_output);

-- MUX_uxn_opcodes_h_l1159_c21_dcf2
MUX_uxn_opcodes_h_l1159_c21_dcf2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1159_c21_dcf2_cond,
MUX_uxn_opcodes_h_l1159_c21_dcf2_iftrue,
MUX_uxn_opcodes_h_l1159_c21_dcf2_iffalse,
MUX_uxn_opcodes_h_l1159_c21_dcf2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade
BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_left,
BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_right,
BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca
result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output,
 n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
 t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output,
 n8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output,
 t8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output,
 n8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_return_output,
 t8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output,
 n8_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output,
 sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_return_output,
 MUX_uxn_opcodes_h_l1159_c21_dcf2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1144_c3_f713 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1148_c3_7589 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1158_c3_df2d : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1162_c3_8eb8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1153_l1150_l1147_l1140_DUPLICATE_b451_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_26fe_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_42d3_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1161_l1153_l1150_l1147_DUPLICATE_cd8d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1153_l1150_DUPLICATE_7a75_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1167_l1136_DUPLICATE_7699_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1162_c3_8eb8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1162_c3_8eb8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1144_c3_f713 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1144_c3_f713;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1148_c3_7589 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1148_c3_7589;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_y := resize(to_signed(-1, 2), 4);
     VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1158_c3_df2d := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1158_c3_df2d;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1153_c11_b258] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_left;
     BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output := BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1153_l1150_DUPLICATE_7a75 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1153_l1150_DUPLICATE_7a75_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1147_c11_c3d5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_left;
     BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output := BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1140_c6_b37c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_left;
     BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output := BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_26fe LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_26fe_return_output := result.is_stack_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_42d3 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_42d3_return_output := result.sp_relative_shift;

     -- sp_relative_shift[uxn_opcodes_h_l1156_c30_890f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_ins;
     sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_x;
     sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_return_output := sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1153_l1150_l1147_l1140_DUPLICATE_b451 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1153_l1150_l1147_l1140_DUPLICATE_b451_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1161_c11_eade] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_left;
     BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output := BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1150_c11_0dd1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1161_l1153_l1150_l1147_DUPLICATE_cd8d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1161_l1153_l1150_l1147_DUPLICATE_cd8d_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1159_c21_06c1] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_left;
     BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_return_output := BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1140_c6_b37c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1147_c11_c3d5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1150_c11_0dd1_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1153_c11_b258_return_output;
     VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1159_c21_06c1_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1161_c11_eade_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_42d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_42d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_42d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_42d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1161_l1153_l1150_l1147_DUPLICATE_cd8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1161_l1153_l1150_l1147_DUPLICATE_cd8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1161_l1153_l1150_l1147_DUPLICATE_cd8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1161_l1153_l1150_l1147_DUPLICATE_cd8d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_26fe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_26fe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_26fe_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1161_l1150_l1147_l1140_DUPLICATE_26fe_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1153_l1150_DUPLICATE_7a75_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1153_l1150_DUPLICATE_7a75_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1153_l1150_l1147_l1140_DUPLICATE_b451_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1153_l1150_l1147_l1140_DUPLICATE_b451_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1153_l1150_l1147_l1140_DUPLICATE_b451_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1153_l1150_l1147_l1140_DUPLICATE_b451_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1156_c30_890f_return_output;
     -- MUX[uxn_opcodes_h_l1159_c21_dcf2] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1159_c21_dcf2_cond <= VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_cond;
     MUX_uxn_opcodes_h_l1159_c21_dcf2_iftrue <= VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_iftrue;
     MUX_uxn_opcodes_h_l1159_c21_dcf2_iffalse <= VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_return_output := MUX_uxn_opcodes_h_l1159_c21_dcf2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1161_c7_49ca] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1153_c7_76c0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1161_c7_49ca] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output;

     -- t8_MUX[uxn_opcodes_h_l1150_c7_a553] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1150_c7_a553_cond <= VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_cond;
     t8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue;
     t8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output := t8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;

     -- n8_MUX[uxn_opcodes_h_l1153_c7_76c0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1153_c7_76c0_cond <= VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_cond;
     n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue;
     n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output := n8_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1161_c7_49ca] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue := VAR_MUX_uxn_opcodes_h_l1159_c21_dcf2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1161_c7_49ca_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1153_c7_76c0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1150_c7_a553] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1153_c7_76c0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1153_c7_76c0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1153_c7_76c0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;

     -- t8_MUX[uxn_opcodes_h_l1147_c7_b81b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond <= VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond;
     t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue;
     t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output := t8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;

     -- n8_MUX[uxn_opcodes_h_l1150_c7_a553] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1150_c7_a553_cond <= VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_cond;
     n8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue;
     n8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output := n8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1153_c7_76c0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1147_c7_b81b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1150_c7_a553] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;

     -- t8_MUX[uxn_opcodes_h_l1140_c2_aa8c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond <= VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond;
     t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue;
     t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output := t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1150_c7_a553] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_return_output := result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;

     -- n8_MUX[uxn_opcodes_h_l1147_c7_b81b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_cond;
     n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue;
     n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output := n8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1150_c7_a553] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1150_c7_a553] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1150_c7_a553_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1140_c2_aa8c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;

     -- n8_MUX[uxn_opcodes_h_l1140_c2_aa8c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond;
     n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue;
     n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output := n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1147_c7_b81b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1147_c7_b81b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1147_c7_b81b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1147_c7_b81b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1147_c7_b81b_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1140_c2_aa8c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1140_c2_aa8c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1140_c2_aa8c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1140_c2_aa8c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1167_l1136_DUPLICATE_7699 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1167_l1136_DUPLICATE_7699_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1140_c2_aa8c_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1167_l1136_DUPLICATE_7699_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1167_l1136_DUPLICATE_7699_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
