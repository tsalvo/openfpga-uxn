-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity rot_0CLK_b288bfb7 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end rot_0CLK_b288bfb7;
architecture arch of rot_0CLK_b288bfb7 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal l8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_l8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2656_c6_5da9]
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2656_c2_9519]
signal l8_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2656_c2_9519]
signal t8_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2656_c2_9519]
signal n8_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(3 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2656_c2_9519]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2669_c11_e276]
signal BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2669_c7_6ab4]
signal l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2669_c7_6ab4]
signal t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2669_c7_6ab4]
signal n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2669_c7_6ab4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2669_c7_6ab4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2669_c7_6ab4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2669_c7_6ab4]
signal result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2669_c7_6ab4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_849a]
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2672_c7_ad0c]
signal l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2672_c7_ad0c]
signal t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2672_c7_ad0c]
signal n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_ad0c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2672_c7_ad0c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2672_c7_ad0c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_ad0c]
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_ad0c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2676_c11_6411]
signal BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2676_c7_035d]
signal l8_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l2676_c7_035d]
signal n8_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2676_c7_035d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2676_c7_035d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2676_c7_035d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2676_c7_035d]
signal result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2676_c7_035d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2678_c30_121e]
signal sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2683_c11_7912]
signal BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output : unsigned(0 downto 0);

-- l8_MUX[uxn_opcodes_h_l2683_c7_c172]
signal l8_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
signal l8_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : unsigned(7 downto 0);
signal l8_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2683_c7_c172]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2683_c7_c172]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : signed(3 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2683_c7_c172]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2683_c7_c172]
signal result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2689_c11_fff9]
signal BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2689_c7_42b2]
signal result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2689_c7_42b2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output : unsigned(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2689_c7_42b2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_188e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_stack_index_flipped := ref_toks_3;
      base.u8_value := ref_toks_4;
      base.is_opc_done := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.stack_address_sp_offset := ref_toks_8;
      base.is_ram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9
BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_left,
BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_right,
BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output);

-- l8_MUX_uxn_opcodes_h_l2656_c2_9519
l8_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
l8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
l8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
l8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- t8_MUX_uxn_opcodes_h_l2656_c2_9519
t8_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
t8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
t8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
t8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- n8_MUX_uxn_opcodes_h_l2656_c2_9519
n8_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
n8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
n8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
n8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519
result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519
result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519
result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519
result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276
BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_left,
BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_right,
BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output);

-- l8_MUX_uxn_opcodes_h_l2669_c7_6ab4
l8_MUX_uxn_opcodes_h_l2669_c7_6ab4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond,
l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue,
l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse,
l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output);

-- t8_MUX_uxn_opcodes_h_l2669_c7_6ab4
t8_MUX_uxn_opcodes_h_l2669_c7_6ab4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond,
t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue,
t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse,
t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output);

-- n8_MUX_uxn_opcodes_h_l2669_c7_6ab4
n8_MUX_uxn_opcodes_h_l2669_c7_6ab4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond,
n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue,
n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse,
n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4
result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4
result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4
result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond,
result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4
result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_left,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_right,
BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output);

-- l8_MUX_uxn_opcodes_h_l2672_c7_ad0c
l8_MUX_uxn_opcodes_h_l2672_c7_ad0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond,
l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue,
l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse,
l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output);

-- t8_MUX_uxn_opcodes_h_l2672_c7_ad0c
t8_MUX_uxn_opcodes_h_l2672_c7_ad0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond,
t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue,
t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse,
t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output);

-- n8_MUX_uxn_opcodes_h_l2672_c7_ad0c
n8_MUX_uxn_opcodes_h_l2672_c7_ad0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond,
n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue,
n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse,
n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c
result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411
BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_left,
BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_right,
BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output);

-- l8_MUX_uxn_opcodes_h_l2676_c7_035d
l8_MUX_uxn_opcodes_h_l2676_c7_035d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2676_c7_035d_cond,
l8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue,
l8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse,
l8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output);

-- n8_MUX_uxn_opcodes_h_l2676_c7_035d
n8_MUX_uxn_opcodes_h_l2676_c7_035d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2676_c7_035d_cond,
n8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue,
n8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse,
n8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d
result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d
result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d
result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2678_c30_121e
sp_relative_shift_uxn_opcodes_h_l2678_c30_121e : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_ins,
sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_x,
sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_y,
sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912
BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_left,
BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_right,
BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output);

-- l8_MUX_uxn_opcodes_h_l2683_c7_c172
l8_MUX_uxn_opcodes_h_l2683_c7_c172 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
l8_MUX_uxn_opcodes_h_l2683_c7_c172_cond,
l8_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue,
l8_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse,
l8_MUX_uxn_opcodes_h_l2683_c7_c172_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172
result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172
result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172
result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_cond,
result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9
BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_left,
BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_right,
BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2
result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_cond,
result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2
result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 l8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output,
 l8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 t8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 n8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output,
 l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output,
 t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output,
 n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output,
 l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output,
 t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output,
 n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output,
 l8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output,
 n8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_return_output,
 sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output,
 l8_MUX_uxn_opcodes_h_l2683_c7_c172_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2661_c3_43c3 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2666_c3_135c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_b9b6 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_8438 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2680_c3_4861 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output : unsigned(0 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : unsigned(7 downto 0);
 variable VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2685_c3_f5cd : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2686_c3_bc2c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2690_c3_0d2c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2689_c7_42b2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2672_l2689_l2656_l2669_DUPLICATE_5d54_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2672_l2669_l2683_DUPLICATE_5379_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2672_l2676_l2669_DUPLICATE_2934_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2689_l2683_l2676_l2672_l2669_DUPLICATE_70a7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2695_l2652_DUPLICATE_dca0_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_l8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_l8 := l8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2680_c3_4861 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2680_c3_4861;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_8438 := resize(to_unsigned(3, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2673_c3_8438;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_right := to_unsigned(5, 3);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_x := signed(std_logic_vector(resize(to_unsigned(3, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_b9b6 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2670_c3_b9b6;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2666_c3_135c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2666_c3_135c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2686_c3_bc2c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2686_c3_bc2c;
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2661_c3_43c3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2661_c3_43c3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_right := to_unsigned(2, 2);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2685_c3_f5cd := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2685_c3_f5cd;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2690_c3_0d2c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2690_c3_0d2c;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_y := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_ins := VAR_ins;
     VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue := l8;
     VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse := l8;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_left := VAR_phase;
     VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue := VAR_previous_stack_read;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2683_c11_7912] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_left;
     BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output := BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2656_c2_9519_return_output := result.is_vram_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2656_c2_9519_return_output := result.is_ram_write;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2672_l2669_l2683_DUPLICATE_5379 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2672_l2669_l2683_DUPLICATE_5379_return_output := result.sp_relative_shift;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2656_c2_9519_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2672_l2676_l2669_DUPLICATE_2934 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2672_l2676_l2669_DUPLICATE_2934_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2676_c11_6411] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_left;
     BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output := BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2689_c7_42b2] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2689_c7_42b2_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2689_c11_fff9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2672_c11_849a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_left;
     BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output := BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2656_c2_9519_return_output := result.is_stack_index_flipped;

     -- sp_relative_shift[uxn_opcodes_h_l2678_c30_121e] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_ins;
     sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_x;
     sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_return_output := sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2656_c6_5da9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_left;
     BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output := BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2672_l2689_l2656_l2669_DUPLICATE_5d54 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2672_l2689_l2656_l2669_DUPLICATE_5d54_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2689_l2683_l2676_l2672_l2669_DUPLICATE_70a7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2689_l2683_l2676_l2672_l2669_DUPLICATE_70a7_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2669_c11_e276] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_left;
     BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output := BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;

     -- Submodule level 1
     VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2656_c6_5da9_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2669_c11_e276_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2672_c11_849a_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2676_c11_6411_return_output;
     VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2683_c11_7912_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2689_c11_fff9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2672_l2669_l2683_DUPLICATE_5379_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2672_l2669_l2683_DUPLICATE_5379_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2672_l2669_l2683_DUPLICATE_5379_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2689_l2683_l2676_l2672_l2669_DUPLICATE_70a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2689_l2683_l2676_l2672_l2669_DUPLICATE_70a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2689_l2683_l2676_l2672_l2669_DUPLICATE_70a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2689_l2683_l2676_l2672_l2669_DUPLICATE_70a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2689_l2683_l2676_l2672_l2669_DUPLICATE_70a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2672_l2676_l2669_DUPLICATE_2934_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2672_l2676_l2669_DUPLICATE_2934_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2672_l2676_l2669_DUPLICATE_2934_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2672_l2689_l2656_l2669_DUPLICATE_5d54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2672_l2689_l2656_l2669_DUPLICATE_5d54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2672_l2689_l2656_l2669_DUPLICATE_5d54_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2672_l2689_l2656_l2669_DUPLICATE_5d54_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2656_c2_9519_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2656_c2_9519_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2656_c2_9519_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2656_c2_9519_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2689_c7_42b2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2678_c30_121e_return_output;
     -- t8_MUX[uxn_opcodes_h_l2672_c7_ad0c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond;
     t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue;
     t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output := t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2689_c7_42b2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2683_c7_c172] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- l8_MUX[uxn_opcodes_h_l2683_c7_c172] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2683_c7_c172_cond <= VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_cond;
     l8_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue;
     l8_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_return_output := l8_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2689_c7_42b2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output;

     -- n8_MUX[uxn_opcodes_h_l2676_c7_035d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2676_c7_035d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_cond;
     n8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue;
     n8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output := n8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2689_c7_42b2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output := result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2676_c7_035d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;

     -- Submodule level 2
     VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2689_c7_42b2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2676_c7_035d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;

     -- l8_MUX[uxn_opcodes_h_l2676_c7_035d] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2676_c7_035d_cond <= VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_cond;
     l8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue;
     l8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output := l8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2672_c7_ad0c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond;
     n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue;
     n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output := n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2683_c7_c172] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_return_output := result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2672_c7_ad0c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;

     -- t8_MUX[uxn_opcodes_h_l2669_c7_6ab4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond <= VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond;
     t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue;
     t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output := t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2683_c7_c172] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2683_c7_c172] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;

     -- Submodule level 3
     VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2683_c7_c172_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2676_c7_035d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2676_c7_035d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;

     -- t8_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     t8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     t8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := t8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2669_c7_6ab4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;

     -- n8_MUX[uxn_opcodes_h_l2669_c7_6ab4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond <= VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond;
     n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue;
     n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output := n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2676_c7_035d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2672_c7_ad0c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;

     -- l8_MUX[uxn_opcodes_h_l2672_c7_ad0c] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond <= VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond;
     l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue;
     l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output := l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;

     -- Submodule level 4
     VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2676_c7_035d_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2672_c7_ad0c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     n8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     n8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := n8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- l8_MUX[uxn_opcodes_h_l2669_c7_6ab4] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond <= VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond;
     l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue;
     l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output := l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2672_c7_ad0c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2672_c7_ad0c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2669_c7_6ab4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;

     -- Submodule level 5
     VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_l8_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2672_c7_ad0c_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2669_c7_6ab4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output := result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2669_c7_6ab4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- l8_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     l8_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     l8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     l8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := l8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2669_c7_6ab4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;

     -- Submodule level 6
     REG_VAR_l8 := VAR_l8_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2669_c7_6ab4_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2656_c2_9519] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_return_output := result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2695_l2652_DUPLICATE_dca0 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2695_l2652_DUPLICATE_dca0_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_188e(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2656_c2_9519_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2656_c2_9519_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2695_l2652_DUPLICATE_dca0_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_188e_uxn_opcodes_h_l2695_l2652_DUPLICATE_dca0_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_l8 <= REG_VAR_l8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     l8 <= REG_COMB_l8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
