-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sth2_0CLK_282a76ca is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end sth2_0CLK_282a76ca;
architecture arch of sth2_0CLK_282a76ca is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2180_c6_f014]
signal BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2180_c2_a34b]
signal t16_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2188_c11_afdc]
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2188_c7_4461]
signal result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2188_c7_4461]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2188_c7_4461]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2188_c7_4461]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2188_c7_4461]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2188_c7_4461]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2188_c7_4461]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2188_c7_4461]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2188_c7_4461]
signal t16_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2190_c30_038b]
signal sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2192_c11_c2ce]
signal BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l2192_c7_45e5]
signal t16_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2200_c11_0654]
signal BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2200_c7_62f0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2200_c7_62f0]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2200_c7_62f0]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2200_c7_62f0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2200_c7_62f0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4a9e( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_sp_shift := ref_toks_6;
      base.is_stack_index_flipped := ref_toks_7;
      base.is_stack_operation_16bit := ref_toks_8;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014
BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_left,
BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_right,
BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b
result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b
result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b
result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b
result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- t16_MUX_uxn_opcodes_h_l2180_c2_a34b
t16_MUX_uxn_opcodes_h_l2180_c2_a34b : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2180_c2_a34b_cond,
t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue,
t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse,
t16_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_left,
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_right,
BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461
result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461
result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- t16_MUX_uxn_opcodes_h_l2188_c7_4461
t16_MUX_uxn_opcodes_h_l2188_c7_4461 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2188_c7_4461_cond,
t16_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue,
t16_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse,
t16_MUX_uxn_opcodes_h_l2188_c7_4461_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2190_c30_038b
sp_relative_shift_uxn_opcodes_h_l2190_c30_038b : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_ins,
sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_x,
sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_y,
sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce
BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_left,
BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_right,
BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5
result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5
result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5
result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5
result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5
result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- t16_MUX_uxn_opcodes_h_l2192_c7_45e5
t16_MUX_uxn_opcodes_h_l2192_c7_45e5 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l2192_c7_45e5_cond,
t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue,
t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse,
t16_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654
BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_left,
BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_right,
BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 t16_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 t16_MUX_uxn_opcodes_h_l2188_c7_4461_return_output,
 sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 t16_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_e8d8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2195_c3_475a : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2197_c3_64f9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2188_l2192_l2180_DUPLICATE_e056_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2192_l2180_DUPLICATE_4b8a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_d86e_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2192_l2180_l2200_DUPLICATE_8b87_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_7f87_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_64ca_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2188_l2192_DUPLICATE_b7c2_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_fdfc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4a9e_uxn_opcodes_h_l2176_l2208_DUPLICATE_3b20_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_right := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_right := to_unsigned(2, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2197_c3_64f9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2197_c3_64f9;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_e8d8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2185_c3_e8d8;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2195_c3_475a := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2195_c3_475a;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_right := to_unsigned(1, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_left := VAR_phase;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := VAR_previous_stack_read;
     VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := t16;
     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2188_l2192_DUPLICATE_b7c2 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2188_l2192_DUPLICATE_b7c2_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l2192_c11_c2ce] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_left;
     BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output := BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2180_c6_f014] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_left;
     BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output := BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_64ca LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_64ca_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2188_c11_afdc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_left;
     BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output := BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2192_l2180_DUPLICATE_4b8a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2192_l2180_DUPLICATE_4b8a_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_7f87 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_7f87_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2188_l2192_l2180_DUPLICATE_e056 LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2188_l2192_l2180_DUPLICATE_e056_return_output := result.u16_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_fdfc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_fdfc_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_d86e LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_d86e_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2200_c11_0654] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_left;
     BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output := BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2190_c30_038b] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_ins;
     sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_x;
     sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_return_output := sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2192_l2180_l2200_DUPLICATE_8b87 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2192_l2180_l2200_DUPLICATE_8b87_return_output := result.is_sp_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2180_c6_f014_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2188_c11_afdc_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2192_c11_c2ce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2200_c11_0654_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2192_l2180_DUPLICATE_4b8a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2192_l2180_DUPLICATE_4b8a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2188_l2192_l2180_DUPLICATE_e056_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2188_l2192_l2180_DUPLICATE_e056_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l2188_l2192_l2180_DUPLICATE_e056_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_64ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_64ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_64ca_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2192_l2180_l2200_DUPLICATE_8b87_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2192_l2180_l2200_DUPLICATE_8b87_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2192_l2180_l2200_DUPLICATE_8b87_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_7f87_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_7f87_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_7f87_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_fdfc_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_fdfc_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l2188_l2192_l2200_DUPLICATE_fdfc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_d86e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_d86e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2188_l2180_l2200_DUPLICATE_d86e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2188_l2192_DUPLICATE_b7c2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2188_l2192_DUPLICATE_b7c2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2190_c30_038b_return_output;
     -- t16_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := t16_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2200_c7_62f0] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2200_c7_62f0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2200_c7_62f0] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2200_c7_62f0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2200_c7_62f0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2200_c7_62f0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- t16_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     t16_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     t16_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := t16_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2192_c7_45e5] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2192_c7_45e5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_t16_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- t16_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := t16_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2188_c7_4461] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2188_c7_4461_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l2180_c2_a34b] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output;

     -- Submodule level 5
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4a9e_uxn_opcodes_h_l2176_l2208_DUPLICATE_3b20 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4a9e_uxn_opcodes_h_l2176_l2208_DUPLICATE_3b20_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4a9e(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l2180_c2_a34b_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4a9e_uxn_opcodes_h_l2176_l2208_DUPLICATE_3b20_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4a9e_uxn_opcodes_h_l2176_l2208_DUPLICATE_3b20_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
