-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity ldz_0CLK_81936ba3 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 previous_ram_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end ldz_0CLK_81936ba3;
architecture arch of ldz_0CLK_81936ba3 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1557_c6_5599]
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1557_c2_9649]
signal tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1557_c2_9649]
signal t8_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1557_c2_9649]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1557_c2_9649]
signal result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1557_c2_9649]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1557_c2_9649]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1557_c2_9649]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1557_c2_9649]
signal result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1557_c2_9649]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1562_c11_16bb]
signal BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal t8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1562_c7_adbb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1565_c11_db4e]
signal BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal t8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : signed(7 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : signed(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1565_c7_6e21]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l1568_c32_e781]
signal BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1568_c32_5919]
signal BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_right : unsigned(0 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1568_c32_8220]
signal MUX_uxn_opcodes_h_l1568_c32_8220_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1568_c32_8220_iftrue : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1568_c32_8220_iffalse : signed(7 downto 0);
signal MUX_uxn_opcodes_h_l1568_c32_8220_return_output : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1571_c11_980b]
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1571_c7_7911]
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1571_c7_7911]
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1571_c7_7911]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1571_c7_7911]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1571_c7_7911]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(0 downto 0);

-- result_ram_addr_MUX[uxn_opcodes_h_l1571_c7_7911]
signal result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(15 downto 0);
signal result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(15 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1571_c7_7911]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1575_c11_1772]
signal BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l1575_c7_19cd]
signal tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(7 downto 0);

-- result_stack_value_MUX[uxn_opcodes_h_l1575_c7_19cd]
signal result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(7 downto 0);
signal result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1575_c7_19cd]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1575_c7_19cd]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(7 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1575_c7_19cd]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1581_c11_17cf]
signal BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1581_c7_12e6]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1581_c7_12e6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output : unsigned(0 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_a287( ref_toks_0 : opcode_result_t;
 ref_toks_1 : signed;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.sp_relative_shift := ref_toks_1;
      base.stack_value := ref_toks_2;
      base.stack_address_sp_offset := ref_toks_3;
      base.is_sp_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.ram_addr := ref_toks_6;
      base.is_opc_done := ref_toks_7;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_left,
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_right,
BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1557_c2_9649
tmp8_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- t8_MUX_uxn_opcodes_h_l1557_c2_9649
t8_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
t8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
t8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
t8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb
BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_left,
BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_right,
BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb
tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- t8_MUX_uxn_opcodes_h_l1562_c7_adbb
t8_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
t8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e
BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_left,
BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_right,
BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21
tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- t8_MUX_uxn_opcodes_h_l1565_c7_6e21
t8_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
t8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781
BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_left,
BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_right,
BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919
BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919 : entity work.BIN_OP_GT_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_left,
BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_right,
BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_return_output);

-- MUX_uxn_opcodes_h_l1568_c32_8220
MUX_uxn_opcodes_h_l1568_c32_8220 : entity work.MUX_uint1_t_int8_t_int8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1568_c32_8220_cond,
MUX_uxn_opcodes_h_l1568_c32_8220_iftrue,
MUX_uxn_opcodes_h_l1568_c32_8220_iffalse,
MUX_uxn_opcodes_h_l1568_c32_8220_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_left,
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_right,
BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1571_c7_7911
tmp8_MUX_uxn_opcodes_h_l1571_c7_7911 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_cond,
tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue,
tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse,
tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_cond,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_return_output);

-- result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_cond,
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue,
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse,
result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772
BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_left,
BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_right,
BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output);

-- tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd
tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_cond,
tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue,
tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse,
tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output);

-- result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_cond,
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue,
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse,
result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf
BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_left,
BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_right,
BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 previous_ram_read,
 -- Registers
 t8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output,
 tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 t8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output,
 tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 t8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output,
 tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 t8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output,
 BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_return_output,
 MUX_uxn_opcodes_h_l1568_c32_8220_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output,
 tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_return_output,
 result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output,
 tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output,
 result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_previous_ram_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_531c : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1563_c3_087b : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : signed(7 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1568_c32_8220_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1568_c32_8220_iftrue : signed(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1568_c32_8220_iffalse : signed(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1568_c32_8220_return_output : signed(7 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_41ec_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(15 downto 0);
 variable VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_cond : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1573_c21_73ee_return_output : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1578_c3_5b94 : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(7 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1557_l1562_l1565_DUPLICATE_6e6a_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1575_DUPLICATE_c893_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_879f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1581_DUPLICATE_4f8c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_f08c_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1581_l1575_DUPLICATE_fb96_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1571_l1575_l1565_DUPLICATE_6018_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a287_uxn_opcodes_h_l1553_l1586_DUPLICATE_9148_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l1568_c32_8220_iffalse := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_right := to_unsigned(3, 2);
     VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_right := to_unsigned(128, 8);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1578_c3_5b94 := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1578_c3_5b94;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_531c := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1559_c3_531c;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1563_c3_087b := resize(to_unsigned(1, 1), 8);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1563_c3_087b;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_right := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1568_c32_8220_iftrue := signed(std_logic_vector(resize(to_unsigned(1, 1), 8)));
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := to_unsigned(1, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;
     VAR_previous_ram_read := previous_ram_read;

     -- Submodule level 0
     VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_left := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_left := VAR_phase;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue := VAR_previous_ram_read;
     VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue := VAR_previous_ram_read;
     VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse := tmp8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1575_DUPLICATE_c893 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1575_DUPLICATE_c893_return_output := result.stack_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_879f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_879f_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1571_c11_980b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1571_l1575_l1565_DUPLICATE_6018 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1571_l1575_l1565_DUPLICATE_6018_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1557_c6_5599] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_left;
     BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output := BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l1568_c32_e781] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_left;
     BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_return_output := BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1565_c11_db4e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_left;
     BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output := BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1581_DUPLICATE_4f8c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1581_DUPLICATE_4f8c_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1581_l1575_DUPLICATE_fb96 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1581_l1575_DUPLICATE_fb96_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1581_c11_17cf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_left;
     BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_return_output := BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1573_c21_73ee] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1573_c21_73ee_return_output := CAST_TO_uint16_t_uint8_t(
     t8);

     -- CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_f08c LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_f08c_return_output := result.ram_addr;

     -- CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1557_l1562_l1565_DUPLICATE_6e6a LATENCY=0
     VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1557_l1562_l1565_DUPLICATE_6e6a_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1562_c11_16bb] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_left;
     BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output := BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1575_c11_1772] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_left;
     BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output := BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output;

     -- CAST_TO_uint16_t[uxn_opcodes_h_l1569_c21_41ec] LATENCY=0
     VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_41ec_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- Submodule level 1
     VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_left := VAR_BIN_OP_AND_uxn_opcodes_h_l1568_c32_e781_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1557_c6_5599_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1562_c11_16bb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1565_c11_db4e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1571_c11_980b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1575_c11_1772_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1581_c11_17cf_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1569_c21_41ec_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue := VAR_CAST_TO_uint16_t_uxn_opcodes_h_l1573_c21_73ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1557_l1562_l1565_DUPLICATE_6e6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1557_l1562_l1565_DUPLICATE_6e6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := VAR_CONST_REF_RD_int8_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1557_l1562_l1565_DUPLICATE_6e6a_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_f08c_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_f08c_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_ram_addr_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_f08c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1581_l1575_DUPLICATE_fb96_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1581_l1575_DUPLICATE_fb96_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1581_l1575_DUPLICATE_fb96_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1581_l1575_DUPLICATE_fb96_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1581_l1575_DUPLICATE_fb96_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_879f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_879f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1557_l1571_l1562_DUPLICATE_879f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1581_DUPLICATE_4f8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1581_DUPLICATE_4f8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1581_DUPLICATE_4f8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1581_DUPLICATE_4f8c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1581_DUPLICATE_4f8c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1571_l1575_l1565_DUPLICATE_6018_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1571_l1575_l1565_DUPLICATE_6018_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1571_l1575_l1565_DUPLICATE_6018_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1575_DUPLICATE_c893_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1575_DUPLICATE_c893_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1575_DUPLICATE_c893_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1575_DUPLICATE_c893_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_stack_value_d41d_uxn_opcodes_h_l1571_l1565_l1562_l1557_l1575_DUPLICATE_c893_return_output;
     -- t8_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := t8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1581_c7_12e6] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1568_c32_5919] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_left;
     BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_return_output := BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1575_c7_19cd] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_cond;
     tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output := tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1575_c7_19cd] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1575_c7_19cd] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output := result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1581_c7_12e6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1571_c7_7911] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1571_c7_7911] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;

     -- Submodule level 2
     VAR_MUX_uxn_opcodes_h_l1568_c32_8220_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1568_c32_5919_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1581_c7_12e6_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1571_c7_7911] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;

     -- MUX[uxn_opcodes_h_l1568_c32_8220] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1568_c32_8220_cond <= VAR_MUX_uxn_opcodes_h_l1568_c32_8220_cond;
     MUX_uxn_opcodes_h_l1568_c32_8220_iftrue <= VAR_MUX_uxn_opcodes_h_l1568_c32_8220_iftrue;
     MUX_uxn_opcodes_h_l1568_c32_8220_iffalse <= VAR_MUX_uxn_opcodes_h_l1568_c32_8220_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1568_c32_8220_return_output := MUX_uxn_opcodes_h_l1568_c32_8220_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1575_c7_19cd] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1575_c7_19cd] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1571_c7_7911] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_cond;
     tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_return_output := tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;

     -- t8_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := t8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1571_c7_7911] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_return_output := result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;

     -- Submodule level 3
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue := VAR_MUX_uxn_opcodes_h_l1568_c32_8220_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1575_c7_19cd_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- t8_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     t8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     t8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := t8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1571_c7_7911] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1571_c7_7911] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1571_c7_7911_return_output;
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_result_ram_addr_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- result_ram_addr_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1565_c7_6e21] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1565_c7_6e21_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_result_stack_value_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1562_c7_adbb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- result_stack_value_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- Submodule level 6
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1562_c7_adbb_return_output;
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1557_c2_9649] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a287_uxn_opcodes_h_l1553_l1586_DUPLICATE_9148 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a287_uxn_opcodes_h_l1553_l1586_DUPLICATE_9148_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a287(
     result,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
     VAR_result_stack_value_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
     VAR_result_ram_addr_MUX_uxn_opcodes_h_l1557_c2_9649_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1557_c2_9649_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a287_uxn_opcodes_h_l1553_l1586_DUPLICATE_9148_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a287_uxn_opcodes_h_l1553_l1586_DUPLICATE_9148_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
