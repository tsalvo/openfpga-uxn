-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity opc_mul_phased_0CLK_c3dfc98c is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(3 downto 0);
 pc : in unsigned(15 downto 0);
 sp : in unsigned(7 downto 0);
 stack_index : in unsigned(0 downto 0);
 ins : in unsigned(7 downto 0);
 k : in unsigned(7 downto 0);
 return_output : out unsigned(0 downto 0));
end opc_mul_phased_0CLK_c3dfc98c;
architecture arch of opc_mul_phased_0CLK_c3dfc98c is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_result : unsigned(0 downto 0);

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_phased_h_l1071_c6_e55f]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1071_c1_c119]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1074_c7_2a45]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1071_c2_3a4f]
signal t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1071_c2_3a4f]
signal n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1071_c2_3a4f]
signal result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output : unsigned(0 downto 0);

-- set_will_fail[uxn_opcodes_phased_h_l1072_c12_5c81]
signal set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_sp : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_k : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_mul : unsigned(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_add : signed(7 downto 0);
signal set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1074_c11_188c]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1074_c1_9d13]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1077_c7_f396]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1074_c7_2a45]
signal t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1074_c7_2a45]
signal n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1074_c7_2a45]
signal result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output : unsigned(0 downto 0);

-- t_register[uxn_opcodes_phased_h_l1075_c8_ff86]
signal t_register_uxn_opcodes_phased_h_l1075_c8_ff86_CLOCK_ENABLE : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_index : unsigned(0 downto 0);
signal t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_ptr : unsigned(7 downto 0);
signal t_register_uxn_opcodes_phased_h_l1075_c8_ff86_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1077_c11_6f26]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1077_c1_9a66]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1080_c7_a86f]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_phased_h_l1077_c7_f396]
signal t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1077_c7_f396]
signal n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1077_c7_f396]
signal result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1078_c8_3f4b]
signal n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1080_c11_630f]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1080_c1_b408]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1083_c7_4280]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_phased_h_l1080_c7_a86f]
signal n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output : unsigned(7 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1080_c7_a86f]
signal result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output : unsigned(0 downto 0);

-- n_register[uxn_opcodes_phased_h_l1081_c8_be9f]
signal n_register_uxn_opcodes_phased_h_l1081_c8_be9f_CLOCK_ENABLE : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_index : unsigned(0 downto 0);
signal n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_ptr : unsigned(7 downto 0);
signal n_register_uxn_opcodes_phased_h_l1081_c8_be9f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1083_c11_aa81]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1083_c1_ee96]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1086_c7_fba4]
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1083_c7_4280]
signal result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output : unsigned(0 downto 0);

-- set[uxn_opcodes_phased_h_l1084_c3_d839]
signal set_uxn_opcodes_phased_h_l1084_c3_d839_CLOCK_ENABLE : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1084_c3_d839_sp : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1084_c3_d839_stack_index : unsigned(0 downto 0);
signal set_uxn_opcodes_phased_h_l1084_c3_d839_ins : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1084_c3_d839_k : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1084_c3_d839_mul : unsigned(7 downto 0);
signal set_uxn_opcodes_phased_h_l1084_c3_d839_add : signed(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1086_c11_139b]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1086_c1_9d7b]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1086_c7_fba4]
signal result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output : unsigned(0 downto 0);

-- BIN_OP_INFERRED_MULT[uxn_opcodes_phased_h_l1087_c33_1ebf]
signal BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_left : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_right : unsigned(7 downto 0);
signal BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_return_output : unsigned(15 downto 0);

-- put_stack[uxn_opcodes_phased_h_l1087_c3_ede9]
signal put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_CLOCK_ENABLE : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_sp : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_stack_index : unsigned(0 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_offset : unsigned(7 downto 0);
signal put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_value : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_phased_h_l1089_c11_f9d4]
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_left : unsigned(3 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_return_output : unsigned(0 downto 0);

-- result_MUX[uxn_opcodes_phased_h_l1089_c7_6ab7]
signal result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_cond : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iftrue : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iffalse : unsigned(0 downto 0);
signal result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_return_output : unsigned(0 downto 0);


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f
BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f
t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond,
t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f
n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond,
n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f
result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond,
result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue,
result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse,
result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output);

-- set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81
set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81 : entity work.set_will_fail_0CLK_23eb2db7 port map (
clk,
set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_CLOCK_ENABLE,
set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_sp,
set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_k,
set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_mul,
set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_add,
set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c
BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c : entity work.BIN_OP_EQ_uint4_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45
t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond,
t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45
n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond,
n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45
result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond,
result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue,
result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse,
result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output);

-- t_register_uxn_opcodes_phased_h_l1075_c8_ff86
t_register_uxn_opcodes_phased_h_l1075_c8_ff86 : entity work.t_register_0CLK_621d5f60 port map (
clk,
t_register_uxn_opcodes_phased_h_l1075_c8_ff86_CLOCK_ENABLE,
t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_index,
t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_ptr,
t_register_uxn_opcodes_phased_h_l1075_c8_ff86_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26
BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26 : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output);

-- t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396
t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond,
t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue,
t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse,
t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396
n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond,
n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1077_c7_f396
result_MUX_uxn_opcodes_phased_h_l1077_c7_f396 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond,
result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue,
result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse,
result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output);

-- n_register_uxn_opcodes_phased_h_l1078_c8_3f4b
n_register_uxn_opcodes_phased_h_l1078_c8_3f4b : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_index,
n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_ptr,
n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f
BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f : entity work.BIN_OP_EQ_uint4_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output);

-- n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f
n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond,
n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue,
n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse,
n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f
result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond,
result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue,
result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse,
result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output);

-- n_register_uxn_opcodes_phased_h_l1081_c8_be9f
n_register_uxn_opcodes_phased_h_l1081_c8_be9f : entity work.n_register_0CLK_621d5f60 port map (
clk,
n_register_uxn_opcodes_phased_h_l1081_c8_be9f_CLOCK_ENABLE,
n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_index,
n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_ptr,
n_register_uxn_opcodes_phased_h_l1081_c8_be9f_return_output);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81
BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_return_output);

-- FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse,
FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1083_c7_4280
result_MUX_uxn_opcodes_phased_h_l1083_c7_4280 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond,
result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue,
result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse,
result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output);

-- set_uxn_opcodes_phased_h_l1084_c3_d839
set_uxn_opcodes_phased_h_l1084_c3_d839 : entity work.set_0CLK_6f2c5aad port map (
clk,
set_uxn_opcodes_phased_h_l1084_c3_d839_CLOCK_ENABLE,
set_uxn_opcodes_phased_h_l1084_c3_d839_sp,
set_uxn_opcodes_phased_h_l1084_c3_d839_stack_index,
set_uxn_opcodes_phased_h_l1084_c3_d839_ins,
set_uxn_opcodes_phased_h_l1084_c3_d839_k,
set_uxn_opcodes_phased_h_l1084_c3_d839_mul,
set_uxn_opcodes_phased_h_l1084_c3_d839_add);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b
BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4
result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond,
result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue,
result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse,
result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output);

-- BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf
BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf : entity work.BIN_OP_INFERRED_MULT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_left,
BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_right,
BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_return_output);

-- put_stack_uxn_opcodes_phased_h_l1087_c3_ede9
put_stack_uxn_opcodes_phased_h_l1087_c3_ede9 : entity work.put_stack_0CLK_b888155f port map (
clk,
put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_CLOCK_ENABLE,
put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_sp,
put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_stack_index,
put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_offset,
put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_value);

-- BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4
BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4 : entity work.BIN_OP_EQ_uint4_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_left,
BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_right,
BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_return_output);

-- result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7
result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_cond,
result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iftrue,
result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iffalse,
result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 pc,
 sp,
 stack_index,
 ins,
 k,
 -- Registers
 n8,
 t8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output,
 result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output,
 set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output,
 result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output,
 t_register_uxn_opcodes_phased_h_l1075_c8_ff86_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output,
 t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output,
 result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output,
 n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output,
 n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output,
 result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output,
 n_register_uxn_opcodes_phased_h_l1081_c8_be9f_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_return_output,
 FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output,
 result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_return_output,
 result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output,
 BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_return_output,
 BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_return_output,
 result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_phase : unsigned(3 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_sp : unsigned(7 downto 0);
 variable VAR_stack_index : unsigned(0 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_k : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_sp : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_k : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_mul : unsigned(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_add : signed(7 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_index : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_ptr : unsigned(7 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_index : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_ptr : unsigned(7 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_sp : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_stack_index : unsigned(0 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_ins : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_k : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_mul : unsigned(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_add : signed(7 downto 0);
 variable VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_sp : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_stack_index : unsigned(0 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_offset : unsigned(7 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_value : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_return_output : unsigned(15 downto 0);
 variable VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_left : unsigned(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_return_output : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iftrue : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iffalse : unsigned(0 downto 0);
 variable VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_cond : unsigned(0 downto 0);
 -- State registers comb logic variables
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_result : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_n8 := n8;
  REG_VAR_t8 := t8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_right := to_unsigned(4, 3);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iffalse := to_unsigned(0, 1);
     VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_add := resize(to_signed(-1, 2), 8);
     VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iftrue := to_unsigned(1, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_right := to_unsigned(1, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_right := to_unsigned(6, 3);
     VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_offset := resize(to_unsigned(0, 1), 8);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_right := to_unsigned(2, 2);
     VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_mul := resize(to_unsigned(2, 2), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_right := to_unsigned(3, 2);
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iffalse := to_unsigned(0, 1);
     VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_add := resize(to_signed(-1, 2), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_pc := pc;
     VAR_sp := sp;
     VAR_stack_index := stack_index;
     VAR_ins := ins;
     VAR_k := k;

     -- Submodule level 0
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iftrue := VAR_CLOCK_ENABLE;
     VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_ins := VAR_ins;
     VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_k := VAR_k;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_k := VAR_k;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_left := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_left := VAR_phase;
     VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue := result;
     VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iffalse := result;
     VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_ptr := VAR_sp;
     VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_sp := VAR_sp;
     VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_sp := VAR_sp;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_sp := VAR_sp;
     VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_ptr := VAR_sp;
     VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_index := VAR_stack_index;
     VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_index := VAR_stack_index;
     VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_stack_index := VAR_stack_index;
     VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_stack_index := VAR_stack_index;
     VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_index := VAR_stack_index;
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_right := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse := t8;
     -- BIN_OP_INFERRED_MULT[uxn_opcodes_phased_h_l1087_c33_1ebf] LATENCY=0
     -- Inputs
     BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_left <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_left;
     BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_right <= VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_right;
     -- Outputs
     VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_return_output := BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1077_c11_6f26] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1083_c11_aa81] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1089_c11_f9d4] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1071_c6_e55f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1080_c11_630f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1086_c11_139b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_return_output;

     -- BIN_OP_EQ[uxn_opcodes_phased_h_l1074_c11_188c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_left <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_left;
     BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_right <= VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output := BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output;

     -- Submodule level 1
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1071_c6_e55f_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1074_c11_188c_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1077_c11_6f26_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1080_c11_630f_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1083_c11_aa81_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1086_c11_139b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_cond := VAR_BIN_OP_EQ_uxn_opcodes_phased_h_l1089_c11_f9d4_return_output;
     VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_value := resize(VAR_BIN_OP_INFERRED_MULT_uxn_opcodes_phased_h_l1087_c33_1ebf_return_output, 8);
     -- result_MUX[uxn_opcodes_phased_h_l1089_c7_6ab7] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_cond;
     result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_return_output := result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1071_c1_c119] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1074_c7_2a45] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;

     -- Submodule level 2
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;
     VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1071_c1_c119_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1089_c7_6ab7_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l1086_c7_fba4] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond;
     result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output := result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1074_c1_9d13] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_return_output;

     -- set_will_fail[uxn_opcodes_phased_h_l1072_c12_5c81] LATENCY=0
     -- Clock enable
     set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_CLOCK_ENABLE <= VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_CLOCK_ENABLE;
     -- Inputs
     set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_sp <= VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_sp;
     set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_k <= VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_k;
     set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_mul <= VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_mul;
     set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_add <= VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_add;
     -- Outputs
     VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_return_output := set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1077_c7_f396] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;

     -- Submodule level 3
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;
     VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1074_c1_9d13_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue := VAR_set_will_fail_uxn_opcodes_phased_h_l1072_c12_5c81_return_output;
     -- t_register[uxn_opcodes_phased_h_l1075_c8_ff86] LATENCY=0
     -- Clock enable
     t_register_uxn_opcodes_phased_h_l1075_c8_ff86_CLOCK_ENABLE <= VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_CLOCK_ENABLE;
     -- Inputs
     t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_index <= VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_index;
     t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_ptr <= VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_stack_ptr;
     -- Outputs
     VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_return_output := t_register_uxn_opcodes_phased_h_l1075_c8_ff86_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1080_c7_a86f] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1077_c1_9a66] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1083_c7_4280] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond;
     result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output := result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output;

     -- Submodule level 4
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1077_c1_9a66_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue := VAR_t_register_uxn_opcodes_phased_h_l1075_c8_ff86_return_output;
     -- n_register[uxn_opcodes_phased_h_l1078_c8_3f4b] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_index;
     n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_return_output := n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1080_c1_b408] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1083_c7_4280] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1080_c7_a86f] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond;
     result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output := result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output;

     -- Submodule level 5
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c7_4280_return_output;
     VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1080_c1_b408_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1078_c8_3f4b_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output;
     -- n_register[uxn_opcodes_phased_h_l1081_c8_be9f] LATENCY=0
     -- Clock enable
     n_register_uxn_opcodes_phased_h_l1081_c8_be9f_CLOCK_ENABLE <= VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_CLOCK_ENABLE;
     -- Inputs
     n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_index <= VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_index;
     n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_ptr <= VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_stack_ptr;
     -- Outputs
     VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_return_output := n_register_uxn_opcodes_phased_h_l1081_c8_be9f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1083_c1_ee96] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1077_c7_f396] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond;
     t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output := t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;

     -- result_MUX[uxn_opcodes_phased_h_l1077_c7_f396] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond;
     result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output := result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1086_c7_fba4] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_cond;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iftrue;
     FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output := FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output;

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c7_fba4_return_output;
     VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1083_c1_ee96_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue := VAR_n_register_uxn_opcodes_phased_h_l1081_c8_be9f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l1074_c7_2a45] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond;
     result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output := result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1074_c7_2a45] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond;
     t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output := t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_phased_h_l1086_c1_9d7b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_return_output;

     -- n8_MUX[uxn_opcodes_phased_h_l1080_c7_a86f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_cond;
     n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output := n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output;

     -- set[uxn_opcodes_phased_h_l1084_c3_d839] LATENCY=0
     -- Clock enable
     set_uxn_opcodes_phased_h_l1084_c3_d839_CLOCK_ENABLE <= VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_CLOCK_ENABLE;
     -- Inputs
     set_uxn_opcodes_phased_h_l1084_c3_d839_sp <= VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_sp;
     set_uxn_opcodes_phased_h_l1084_c3_d839_stack_index <= VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_stack_index;
     set_uxn_opcodes_phased_h_l1084_c3_d839_ins <= VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_ins;
     set_uxn_opcodes_phased_h_l1084_c3_d839_k <= VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_k;
     set_uxn_opcodes_phased_h_l1084_c3_d839_mul <= VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_mul;
     set_uxn_opcodes_phased_h_l1084_c3_d839_add <= VAR_set_uxn_opcodes_phased_h_l1084_c3_d839_add;
     -- Outputs

     -- Submodule level 7
     VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_phased_h_l1086_c1_9d7b_return_output;
     VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1080_c7_a86f_return_output;
     VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse := VAR_result_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;
     VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse := VAR_t8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;
     -- result_MUX[uxn_opcodes_phased_h_l1071_c2_3a4f] LATENCY=0
     -- Inputs
     result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond <= VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond;
     result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue <= VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue;
     result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse <= VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse;
     -- Outputs
     VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output := result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output;

     -- t8_MUX[uxn_opcodes_phased_h_l1071_c2_3a4f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond <= VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond;
     t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue <= VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue;
     t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse <= VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output := t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output;

     -- put_stack[uxn_opcodes_phased_h_l1087_c3_ede9] LATENCY=0
     -- Clock enable
     put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_CLOCK_ENABLE <= VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_CLOCK_ENABLE;
     -- Inputs
     put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_sp <= VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_sp;
     put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_stack_index <= VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_stack_index;
     put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_offset <= VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_offset;
     put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_value <= VAR_put_stack_uxn_opcodes_phased_h_l1087_c3_ede9_value;
     -- Outputs

     -- n8_MUX[uxn_opcodes_phased_h_l1077_c7_f396] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_cond;
     n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output := n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;

     -- Submodule level 8
     VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1077_c7_f396_return_output;
     REG_VAR_result := VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output;
     VAR_return_output := VAR_result_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1074_c7_2a45] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_cond;
     n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output := n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;

     -- Submodule level 9
     VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse := VAR_n8_MUX_uxn_opcodes_phased_h_l1074_c7_2a45_return_output;
     -- n8_MUX[uxn_opcodes_phased_h_l1071_c2_3a4f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond <= VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_cond;
     n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue <= VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iftrue;
     n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse <= VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output := n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output;

     -- Submodule level 10
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_phased_h_l1071_c2_3a4f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     n8 <= REG_COMB_n8;
     t8 <= REG_COMB_t8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
