-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 35
entity jmp2_0CLK_d6642053 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end jmp2_0CLK_d6642053;
architecture arch of jmp2_0CLK_d6642053 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l645_c6_d898]
signal BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l645_c2_6b81]
signal result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l645_c2_6b81]
signal t16_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l658_c11_0667]
signal BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l658_c7_20c6]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(3 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l658_c7_20c6]
signal result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(15 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l658_c7_20c6]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : signed(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l658_c7_20c6]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l658_c7_20c6]
signal result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l658_c7_20c6]
signal t16_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l661_c11_957d]
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l661_c7_283d]
signal result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l661_c7_283d]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l661_c7_283d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l661_c7_283d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_return_output : signed(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l661_c7_283d]
signal t16_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l661_c7_283d_return_output : unsigned(15 downto 0);

-- CONST_SL_8[uxn_opcodes_h_l663_c3_0ef6]
signal CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_x : unsigned(15 downto 0);
signal CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l665_c11_eafc]
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l665_c7_126c]
signal result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l665_c7_126c]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l665_c7_126c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l665_c7_126c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_return_output : signed(3 downto 0);

-- t16_MUX[uxn_opcodes_h_l665_c7_126c]
signal t16_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l665_c7_126c_return_output : unsigned(15 downto 0);

-- BIN_OP_OR[uxn_opcodes_h_l666_c3_8d4d]
signal BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_left : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_right : unsigned(15 downto 0);
signal BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l667_c30_319a]
signal sp_relative_shift_uxn_opcodes_h_l667_c30_319a_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l667_c30_319a_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l667_c30_319a_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l667_c30_319a_return_output : signed(3 downto 0);

function CAST_TO_uint16_t_uint8_t( rhs : unsigned) return unsigned is

  --variable rhs : unsigned(7 downto 0);
  variable return_output : unsigned(15 downto 0);

begin

      return_output := unsigned(std_logic_vector(resize(rhs,16)));
    return return_output;
end function;

function CONST_REF_RD_opcode_result_t_opcode_result_t_5ddc( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.is_stack_index_flipped := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.u16_value := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898
BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_left,
BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_right,
BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81
result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81
result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81
result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81
result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81
result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81
result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81
result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- t16_MUX_uxn_opcodes_h_l645_c2_6b81
t16_MUX_uxn_opcodes_h_l645_c2_6b81 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l645_c2_6b81_cond,
t16_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue,
t16_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse,
t16_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667
BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_left,
BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_right,
BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6
result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_cond,
result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6
result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6
result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6
result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_return_output);

-- t16_MUX_uxn_opcodes_h_l658_c7_20c6
t16_MUX_uxn_opcodes_h_l658_c7_20c6 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l658_c7_20c6_cond,
t16_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue,
t16_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse,
t16_MUX_uxn_opcodes_h_l658_c7_20c6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d
BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_left,
BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_right,
BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d
result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_cond,
result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_return_output);

-- t16_MUX_uxn_opcodes_h_l661_c7_283d
t16_MUX_uxn_opcodes_h_l661_c7_283d : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l661_c7_283d_cond,
t16_MUX_uxn_opcodes_h_l661_c7_283d_iftrue,
t16_MUX_uxn_opcodes_h_l661_c7_283d_iffalse,
t16_MUX_uxn_opcodes_h_l661_c7_283d_return_output);

-- CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6
CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6 : entity work.CONST_SL_8_uint16_t_0CLK_de264c78 port map (
CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_x,
CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc
BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_left,
BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_right,
BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c
result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_cond,
result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_return_output);

-- t16_MUX_uxn_opcodes_h_l665_c7_126c
t16_MUX_uxn_opcodes_h_l665_c7_126c : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l665_c7_126c_cond,
t16_MUX_uxn_opcodes_h_l665_c7_126c_iftrue,
t16_MUX_uxn_opcodes_h_l665_c7_126c_iffalse,
t16_MUX_uxn_opcodes_h_l665_c7_126c_return_output);

-- BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d
BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d : entity work.BIN_OP_OR_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_left,
BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_right,
BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l667_c30_319a
sp_relative_shift_uxn_opcodes_h_l667_c30_319a : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l667_c30_319a_ins,
sp_relative_shift_uxn_opcodes_h_l667_c30_319a_x,
sp_relative_shift_uxn_opcodes_h_l667_c30_319a_y,
sp_relative_shift_uxn_opcodes_h_l667_c30_319a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 t16_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_return_output,
 t16_MUX_uxn_opcodes_h_l658_c7_20c6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_return_output,
 t16_MUX_uxn_opcodes_h_l661_c7_283d_return_output,
 CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_return_output,
 t16_MUX_uxn_opcodes_h_l665_c7_126c_return_output,
 BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_return_output,
 sp_relative_shift_uxn_opcodes_h_l667_c30_319a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l650_c3_e507 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l655_c3_b30e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l659_c3_b786 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l658_c7_20c6_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_cond : unsigned(0 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_return_output : unsigned(15 downto 0);
 variable VAR_CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_x : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_return_output : unsigned(15 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l661_l645_l665_l658_DUPLICATE_9a9a_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_382a_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_963c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_83b9_return_output : unsigned(0 downto 0);
 variable VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l662_l666_DUPLICATE_8db0_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5ddc_uxn_opcodes_h_l641_l673_DUPLICATE_9c8a_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l655_c3_b30e := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l655_c3_b30e;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iftrue := to_unsigned(1, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l650_c3_e507 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l650_c3_e507;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l659_c3_b786 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l659_c3_b786;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_y := resize(to_signed(-2, 3), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_ins := VAR_ins;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_left := VAR_phase;
     VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_left := t16;
     VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_iffalse := t16;
     -- BIN_OP_EQ[uxn_opcodes_h_l665_c11_eafc] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_left;
     BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output := BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l661_l645_l665_l658_DUPLICATE_9a9a LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l661_l645_l665_l658_DUPLICATE_9a9a_return_output := result.u16_value;

     -- result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output := result.is_stack_write;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l645_c2_6b81_return_output := result.is_stack_index_flipped;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_83b9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_83b9_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_963c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_963c_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l667_c30_319a] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l667_c30_319a_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_ins;
     sp_relative_shift_uxn_opcodes_h_l667_c30_319a_x <= VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_x;
     sp_relative_shift_uxn_opcodes_h_l667_c30_319a_y <= VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_return_output := sp_relative_shift_uxn_opcodes_h_l667_c30_319a_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l658_c11_0667] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_left;
     BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output := BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output;

     -- CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l662_l666_DUPLICATE_8db0 LATENCY=0
     VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l662_l666_DUPLICATE_8db0_return_output := CAST_TO_uint16_t_uint8_t(
     VAR_previous_stack_read);

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l658_c7_20c6] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l658_c7_20c6_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l661_c11_957d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_left;
     BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output := BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l645_c6_d898] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_left;
     BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output := BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_382a LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_382a_return_output := result.sp_relative_shift;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l645_c6_d898_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l658_c11_0667_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l661_c11_957d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l665_c11_eafc_return_output;
     VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_right := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l662_l666_DUPLICATE_8db0_return_output;
     VAR_CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_x := VAR_CAST_TO_uint16_t_uint8_t_uxn_opcodes_h_l662_l666_DUPLICATE_8db0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_382a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_382a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_382a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l661_l645_l665_l658_DUPLICATE_9a9a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l661_l645_l665_l658_DUPLICATE_9a9a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l661_l645_l665_l658_DUPLICATE_9a9a_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l661_l645_l665_l658_DUPLICATE_9a9a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_83b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_83b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_83b9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_963c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_963c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l661_l665_l658_DUPLICATE_963c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l645_c2_6b81_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_is_stack_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l645_c2_6b81_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l658_c7_20c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l667_c30_319a_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l665_c7_126c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l665_c7_126c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l665_c7_126c] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_return_output;

     -- CONST_SL_8[uxn_opcodes_h_l663_c3_0ef6] LATENCY=0
     -- Inputs
     CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_x <= VAR_CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_x;
     -- Outputs
     VAR_CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_return_output := CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- BIN_OP_OR[uxn_opcodes_h_l666_c3_8d4d] LATENCY=0
     -- Inputs
     BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_left <= VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_left;
     BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_right <= VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_right;
     -- Outputs
     VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_return_output := BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l658_c7_20c6] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;

     -- Submodule level 2
     VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_iftrue := VAR_BIN_OP_OR_uxn_opcodes_h_l666_c3_8d4d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_iftrue := VAR_CONST_SL_8_uxn_opcodes_h_l663_c3_0ef6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l665_c7_126c_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l665_c7_126c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l665_c7_126c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l661_c7_283d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l661_c7_283d] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_return_output;

     -- t16_MUX[uxn_opcodes_h_l665_c7_126c] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l665_c7_126c_cond <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_cond;
     t16_MUX_uxn_opcodes_h_l665_c7_126c_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_iftrue;
     t16_MUX_uxn_opcodes_h_l665_c7_126c_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_return_output := t16_MUX_uxn_opcodes_h_l665_c7_126c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l665_c7_126c] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_cond;
     result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_return_output := result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l661_c7_283d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l661_c7_283d_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l661_c7_283d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l661_c7_283d_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l665_c7_126c_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_iffalse := VAR_t16_MUX_uxn_opcodes_h_l665_c7_126c_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l658_c7_20c6] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l661_c7_283d] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_cond;
     result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_return_output := result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l658_c7_20c6] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;

     -- t16_MUX[uxn_opcodes_h_l661_c7_283d] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l661_c7_283d_cond <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_cond;
     t16_MUX_uxn_opcodes_h_l661_c7_283d_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_iftrue;
     t16_MUX_uxn_opcodes_h_l661_c7_283d_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_return_output := t16_MUX_uxn_opcodes_h_l661_c7_283d_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l658_c7_20c6] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l661_c7_283d_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse := VAR_t16_MUX_uxn_opcodes_h_l661_c7_283d_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l658_c7_20c6] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_cond;
     result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_return_output := result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- t16_MUX[uxn_opcodes_h_l658_c7_20c6] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l658_c7_20c6_cond <= VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_cond;
     t16_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_iftrue;
     t16_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_return_output := t16_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;

     -- Submodule level 5
     VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse := VAR_t16_MUX_uxn_opcodes_h_l658_c7_20c6_return_output;
     -- t16_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     t16_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     t16_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := t16_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l645_c2_6b81] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_cond;
     result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_return_output := result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;

     -- Submodule level 6
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l645_c2_6b81_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5ddc_uxn_opcodes_h_l641_l673_DUPLICATE_9c8a LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5ddc_uxn_opcodes_h_l641_l673_DUPLICATE_9c8a_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5ddc(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l645_c2_6b81_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l645_c2_6b81_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5ddc_uxn_opcodes_h_l641_l673_DUPLICATE_9c8a_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5ddc_uxn_opcodes_h_l641_l673_DUPLICATE_9c8a_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
