-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 50
entity and_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_fedec265;
architecture arch of and_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l950_c6_51fd]
signal BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l950_c2_f139]
signal n8_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l950_c2_f139]
signal t8_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l950_c2_f139]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l950_c2_f139]
signal result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l950_c2_f139]
signal result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l950_c2_f139]
signal result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l950_c2_f139]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l950_c2_f139]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l955_c11_74e3]
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l955_c7_b890]
signal n8_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l955_c7_b890]
signal t8_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l955_c7_b890]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l955_c7_b890]
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l955_c7_b890]
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l955_c7_b890]
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l955_c7_b890]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l955_c7_b890]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l958_c11_74a7]
signal BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l958_c7_fcdf]
signal n8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l958_c7_fcdf]
signal t8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l958_c7_fcdf]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l958_c7_fcdf]
signal result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l958_c7_fcdf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l958_c7_fcdf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l958_c7_fcdf]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l958_c7_fcdf]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l962_c11_ba19]
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l962_c7_3a6a]
signal n8_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l962_c7_3a6a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l962_c7_3a6a]
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l962_c7_3a6a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l962_c7_3a6a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l962_c7_3a6a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l962_c7_3a6a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l965_c11_698d]
signal BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l965_c7_fd36]
signal n8_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l965_c7_fd36]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l965_c7_fd36]
signal result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l965_c7_fd36]
signal result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l965_c7_fd36]
signal result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l965_c7_fd36]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l965_c7_fd36]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l968_c30_94dc]
signal sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l971_c21_f8a9]
signal BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l973_c11_ae39]
signal BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l973_c7_beaf]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l973_c7_beaf]
signal result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l973_c7_beaf]
signal result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd
BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_left,
BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_right,
BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output);

-- n8_MUX_uxn_opcodes_h_l950_c2_f139
n8_MUX_uxn_opcodes_h_l950_c2_f139 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l950_c2_f139_cond,
n8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue,
n8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse,
n8_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

-- t8_MUX_uxn_opcodes_h_l950_c2_f139
t8_MUX_uxn_opcodes_h_l950_c2_f139 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l950_c2_f139_cond,
t8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue,
t8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse,
t8_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139
result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_cond,
result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139
result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139
result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139
result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139
result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3
BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_left,
BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_right,
BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output);

-- n8_MUX_uxn_opcodes_h_l955_c7_b890
n8_MUX_uxn_opcodes_h_l955_c7_b890 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l955_c7_b890_cond,
n8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue,
n8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse,
n8_MUX_uxn_opcodes_h_l955_c7_b890_return_output);

-- t8_MUX_uxn_opcodes_h_l955_c7_b890
t8_MUX_uxn_opcodes_h_l955_c7_b890 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l955_c7_b890_cond,
t8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue,
t8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse,
t8_MUX_uxn_opcodes_h_l955_c7_b890_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890
result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_cond,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7
BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_left,
BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_right,
BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output);

-- n8_MUX_uxn_opcodes_h_l958_c7_fcdf
n8_MUX_uxn_opcodes_h_l958_c7_fcdf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond,
n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue,
n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse,
n8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output);

-- t8_MUX_uxn_opcodes_h_l958_c7_fcdf
t8_MUX_uxn_opcodes_h_l958_c7_fcdf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond,
t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue,
t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse,
t8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf
result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_cond,
result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf
result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf
result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf
result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf
result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19
BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_left,
BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_right,
BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output);

-- n8_MUX_uxn_opcodes_h_l962_c7_3a6a
n8_MUX_uxn_opcodes_h_l962_c7_3a6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l962_c7_3a6a_cond,
n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue,
n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse,
n8_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a
result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_cond,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d
BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_left,
BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_right,
BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output);

-- n8_MUX_uxn_opcodes_h_l965_c7_fd36
n8_MUX_uxn_opcodes_h_l965_c7_fd36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l965_c7_fd36_cond,
n8_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue,
n8_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse,
n8_MUX_uxn_opcodes_h_l965_c7_fd36_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36
result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_cond,
result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36
result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36
result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36
result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36
result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output);

-- sp_relative_shift_uxn_opcodes_h_l968_c30_94dc
sp_relative_shift_uxn_opcodes_h_l968_c30_94dc : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_ins,
sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_x,
sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_y,
sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9
BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9 : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_left,
BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_right,
BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39
BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_left,
BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_right,
BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf
result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf
result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf
result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output,
 n8_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
 t8_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output,
 n8_MUX_uxn_opcodes_h_l955_c7_b890_return_output,
 t8_MUX_uxn_opcodes_h_l955_c7_b890_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output,
 n8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output,
 t8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output,
 n8_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output,
 n8_MUX_uxn_opcodes_h_l965_c7_fd36_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output,
 sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_return_output,
 BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l952_c3_1720 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l956_c3_f9d5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_3bfa : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l963_c3_bfe0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l970_c3_f6c3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l965_c7_fd36_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_5b43_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_1d30_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_b815_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_4731_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l965_l962_l958_l955_l973_DUPLICATE_f73a_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l979_l946_DUPLICATE_d79d_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_right := to_unsigned(5, 3);
     VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_right := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l952_c3_1720 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l952_c3_1720;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l970_c3_f6c3 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l970_c3_f6c3;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_3bfa := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l960_c3_3bfa;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l956_c3_f9d5 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l956_c3_f9d5;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l963_c3_bfe0 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l963_c3_bfe0;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l965_l962_l958_l955_l973_DUPLICATE_f73a LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l965_l962_l958_l955_l973_DUPLICATE_f73a_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_5b43 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_5b43_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_1d30 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_1d30_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l958_c11_74a7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_left;
     BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output := BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l965_c7_fd36] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l965_c7_fd36_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l955_c11_74e3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_left;
     BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output := BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l973_c11_ae39] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_left;
     BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output := BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_b815 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_b815_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_4731 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_4731_return_output := result.is_sp_shift;

     -- sp_relative_shift[uxn_opcodes_h_l968_c30_94dc] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_ins;
     sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_x <= VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_x;
     sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_y <= VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_return_output := sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l962_c11_ba19] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_left;
     BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output := BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output;

     -- BIN_OP_AND[uxn_opcodes_h_l971_c21_f8a9] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_left;
     BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_return_output := BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l950_c6_51fd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_left;
     BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output := BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l965_c11_698d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_left;
     BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output := BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l971_c21_f8a9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l950_c6_51fd_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l955_c11_74e3_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l958_c11_74a7_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l962_c11_ba19_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l965_c11_698d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l973_c11_ae39_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_b815_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_b815_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_b815_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_b815_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_b815_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l965_l962_l958_l955_l973_DUPLICATE_f73a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l965_l962_l958_l955_l973_DUPLICATE_f73a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l965_l962_l958_l955_l973_DUPLICATE_f73a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l965_l962_l958_l955_l973_DUPLICATE_f73a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l965_l962_l958_l955_l973_DUPLICATE_f73a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_4731_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_4731_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_4731_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_4731_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_4731_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_1d30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_1d30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_1d30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_1d30_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l962_l958_l955_l950_l973_DUPLICATE_1d30_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_5b43_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_5b43_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_5b43_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_5b43_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l965_l962_l958_l955_l950_DUPLICATE_5b43_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l965_c7_fd36_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l968_c30_94dc_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l965_c7_fd36] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l973_c7_beaf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l965_c7_fd36] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l965_c7_fd36] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_cond;
     result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_return_output := result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l973_c7_beaf] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_return_output;

     -- t8_MUX[uxn_opcodes_h_l958_c7_fcdf] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond <= VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond;
     t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue;
     t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output := t8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l973_c7_beaf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_return_output;

     -- n8_MUX[uxn_opcodes_h_l965_c7_fd36] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l965_c7_fd36_cond <= VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_cond;
     n8_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue;
     n8_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_return_output := n8_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l973_c7_beaf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l973_c7_beaf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l973_c7_beaf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse := VAR_t8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l962_c7_3a6a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l962_c7_3a6a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;

     -- n8_MUX[uxn_opcodes_h_l962_c7_3a6a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l962_c7_3a6a_cond <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_cond;
     n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue;
     n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output := n8_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l965_c7_fd36] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l965_c7_fd36] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;

     -- t8_MUX[uxn_opcodes_h_l955_c7_b890] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l955_c7_b890_cond <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_cond;
     t8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue;
     t8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_return_output := t8_MUX_uxn_opcodes_h_l955_c7_b890_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l962_c7_3a6a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output := result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l965_c7_fd36] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse := VAR_n8_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l965_c7_fd36_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse := VAR_t8_MUX_uxn_opcodes_h_l955_c7_b890_return_output;
     -- n8_MUX[uxn_opcodes_h_l958_c7_fcdf] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond <= VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_cond;
     n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue;
     n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output := n8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l962_c7_3a6a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l962_c7_3a6a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;

     -- t8_MUX[uxn_opcodes_h_l950_c2_f139] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l950_c2_f139_cond <= VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_cond;
     t8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue;
     t8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_return_output := t8_MUX_uxn_opcodes_h_l950_c2_f139_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l958_c7_fcdf] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l958_c7_fcdf] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l962_c7_3a6a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l958_c7_fcdf] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_cond;
     result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output := result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse := VAR_n8_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l962_c7_3a6a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l950_c2_f139_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l955_c7_b890] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l958_c7_fcdf] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l958_c7_fcdf] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l955_c7_b890] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_cond;
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_return_output := result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l958_c7_fcdf] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l955_c7_b890] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output;

     -- n8_MUX[uxn_opcodes_h_l955_c7_b890] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l955_c7_b890_cond <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_cond;
     n8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_iftrue;
     n8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_return_output := n8_MUX_uxn_opcodes_h_l955_c7_b890_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse := VAR_n8_MUX_uxn_opcodes_h_l955_c7_b890_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l958_c7_fcdf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l955_c7_b890_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l955_c7_b890_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l950_c2_f139] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l955_c7_b890] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l950_c2_f139] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l955_c7_b890] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l950_c2_f139] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_cond;
     result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_return_output := result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_return_output;

     -- n8_MUX[uxn_opcodes_h_l950_c2_f139] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l950_c2_f139_cond <= VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_cond;
     n8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_iftrue;
     n8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_return_output := n8_MUX_uxn_opcodes_h_l950_c2_f139_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l955_c7_b890] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l950_c2_f139_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l955_c7_b890_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l955_c7_b890_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l955_c7_b890_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l950_c2_f139] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l950_c2_f139] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l950_c2_f139] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l979_l946_DUPLICATE_d79d LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l979_l946_DUPLICATE_d79d_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l950_c2_f139_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l979_l946_DUPLICATE_d79d_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l979_l946_DUPLICATE_d79d_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
