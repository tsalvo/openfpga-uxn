-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity sft_0CLK_46cced44 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sft_0CLK_46cced44;
architecture arch of sft_0CLK_46cced44 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal tmp8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_tmp8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2236_c6_5798]
signal BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : signed(3 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(7 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(3 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2236_c2_5e7c]
signal tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2249_c11_04f8]
signal BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2249_c7_1432]
signal n8_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2249_c7_1432]
signal t8_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2249_c7_1432]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2249_c7_1432]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2249_c7_1432]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2249_c7_1432]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2249_c7_1432]
signal result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2249_c7_1432]
signal tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2252_c11_4d69]
signal BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2252_c7_c2ab]
signal n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2252_c7_c2ab]
signal t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2252_c7_c2ab]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2252_c7_c2ab]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2252_c7_c2ab]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2252_c7_c2ab]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2252_c7_c2ab]
signal result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2252_c7_c2ab]
signal tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2254_c30_c3c4]
signal sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2256_c11_d531]
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2256_c7_e6a8]
signal n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2256_c7_e6a8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2256_c7_e6a8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2256_c7_e6a8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : signed(3 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2256_c7_e6a8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2256_c7_e6a8]
signal result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(7 downto 0);

-- tmp8_MUX[uxn_opcodes_h_l2256_c7_e6a8]
signal tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(7 downto 0);
signal tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(7 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l2259_c18_a8de]
signal BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_return_output : unsigned(7 downto 0);

-- BIN_OP_SR[uxn_opcodes_h_l2259_c11_1037]
signal BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_left : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_right : unsigned(7 downto 0);
signal BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_return_output : unsigned(7 downto 0);

-- CONST_SR_4[uxn_opcodes_h_l2259_c34_d847]
signal CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_x : unsigned(7 downto 0);
signal CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_return_output : unsigned(7 downto 0);

-- BIN_OP_SL[uxn_opcodes_h_l2259_c11_4f50]
signal BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_left : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_right : unsigned(7 downto 0);
signal BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_e848( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.is_ram_write := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_vram_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.is_stack_index_flipped := ref_toks_6;
      base.stack_address_sp_offset := ref_toks_7;
      base.is_pc_updated := ref_toks_8;
      base.is_opc_done := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798
BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_left,
BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_right,
BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output);

-- n8_MUX_uxn_opcodes_h_l2236_c2_5e7c
n8_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- t8_MUX_uxn_opcodes_h_l2236_c2_5e7c
t8_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c
tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond,
tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue,
tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse,
tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8
BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_left,
BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_right,
BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output);

-- n8_MUX_uxn_opcodes_h_l2249_c7_1432
n8_MUX_uxn_opcodes_h_l2249_c7_1432 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2249_c7_1432_cond,
n8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue,
n8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse,
n8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output);

-- t8_MUX_uxn_opcodes_h_l2249_c7_1432
t8_MUX_uxn_opcodes_h_l2249_c7_1432 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2249_c7_1432_cond,
t8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue,
t8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse,
t8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_cond,
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2249_c7_1432
tmp8_MUX_uxn_opcodes_h_l2249_c7_1432 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_cond,
tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue,
tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse,
tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69
BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_left,
BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_right,
BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output);

-- n8_MUX_uxn_opcodes_h_l2252_c7_c2ab
n8_MUX_uxn_opcodes_h_l2252_c7_c2ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond,
n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue,
n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse,
n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output);

-- t8_MUX_uxn_opcodes_h_l2252_c7_c2ab
t8_MUX_uxn_opcodes_h_l2252_c7_c2ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond,
t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue,
t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse,
t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond,
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab
tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond,
tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue,
tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse,
tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4
sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_ins,
sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_x,
sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_y,
sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_left,
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_right,
BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output);

-- n8_MUX_uxn_opcodes_h_l2256_c7_e6a8
n8_MUX_uxn_opcodes_h_l2256_c7_e6a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond,
n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue,
n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse,
n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond,
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output);

-- tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8
tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond,
tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue,
tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse,
tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de
BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_left,
BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_right,
BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_return_output);

-- BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037
BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037 : entity work.BIN_OP_SR_uint8_t_uint8_t_0CLK_25d197a7 port map (
BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_left,
BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_right,
BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_return_output);

-- CONST_SR_4_uxn_opcodes_h_l2259_c34_d847
CONST_SR_4_uxn_opcodes_h_l2259_c34_d847 : entity work.CONST_SR_4_uint8_t_0CLK_de264c78 port map (
CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_x,
CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_return_output);

-- BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50
BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50 : entity work.BIN_OP_SL_uint8_t_uint8_t_0CLK_10d8c973 port map (
BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_left,
BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_right,
BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 tmp8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output,
 n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output,
 n8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output,
 t8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_return_output,
 tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output,
 n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output,
 t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output,
 tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output,
 sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output,
 n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output,
 tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output,
 BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_return_output,
 BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_return_output,
 CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_return_output,
 BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2241_c3_01e8 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2246_c3_0d85 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2250_c3_a21f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_7169 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2258_c3_088b : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse : unsigned(7 downto 0);
 variable VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_left : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_right : unsigned(7 downto 0);
 variable VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_x : unsigned(7 downto 0);
 variable VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2252_l2236_l2256_l2249_DUPLICATE_48a0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_1d83_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_7fe4_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_02e7_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2252_l2256_DUPLICATE_d4e0_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2232_l2266_DUPLICATE_340f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_tmp8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_tmp8 := tmp8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2241_c3_01e8 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2241_c3_01e8;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_right := to_unsigned(15, 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := to_unsigned(0, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2250_c3_a21f := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2250_c3_a21f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2246_c3_0d85 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2246_c3_0d85;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_7169 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2261_c3_7169;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_right := to_unsigned(2, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2258_c3_088b := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2258_c3_088b;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_left := VAR_phase;
     VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_left := t8;
     VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_x := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse := t8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue := tmp8;
     VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse := tmp8;
     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2252_l2236_l2256_l2249_DUPLICATE_48a0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2252_l2236_l2256_l2249_DUPLICATE_48a0_return_output := result.u8_value;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_1d83 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_1d83_return_output := result.is_stack_write;

     -- sp_relative_shift[uxn_opcodes_h_l2254_c30_c3c4] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_ins;
     sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_x;
     sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_return_output := sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2249_c11_04f8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_left;
     BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output := BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_7fe4 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_7fe4_return_output := result.sp_relative_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l2259_c18_a8de] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_left;
     BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_return_output := BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2252_l2256_DUPLICATE_d4e0 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2252_l2256_DUPLICATE_d4e0_return_output := result.stack_address_sp_offset;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output := result.is_vram_write;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output := result.is_ram_write;

     -- CONST_SR_4[uxn_opcodes_h_l2259_c34_d847] LATENCY=0
     -- Inputs
     CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_x <= VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_x;
     -- Outputs
     VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_return_output := CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_02e7 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_02e7_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l2256_c11_d531] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_left;
     BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output := BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2252_c11_4d69] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_left;
     BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output := BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2236_c6_5798] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_left;
     BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output := BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;

     -- Submodule level 1
     VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_right := VAR_BIN_OP_AND_uxn_opcodes_h_l2259_c18_a8de_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2236_c6_5798_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2249_c11_04f8_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2252_c11_4d69_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2256_c11_d531_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_7fe4_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2256_l2249_DUPLICATE_7fe4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_02e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_02e7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_02e7_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_1d83_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_1d83_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2252_l2256_l2249_DUPLICATE_1d83_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2252_l2256_DUPLICATE_d4e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2252_l2256_DUPLICATE_d4e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2252_l2236_l2256_l2249_DUPLICATE_48a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2252_l2236_l2256_l2249_DUPLICATE_48a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2252_l2236_l2256_l2249_DUPLICATE_48a0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2252_l2236_l2256_l2249_DUPLICATE_48a0_return_output;
     VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_right := VAR_CONST_SR_4_uxn_opcodes_h_l2259_c34_d847_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2236_c2_5e7c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2254_c30_c3c4_return_output;
     -- BIN_OP_SR[uxn_opcodes_h_l2259_c11_1037] LATENCY=0
     -- Inputs
     BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_left <= VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_left;
     BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_right <= VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_right;
     -- Outputs
     VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_return_output := BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_return_output;

     -- t8_MUX[uxn_opcodes_h_l2252_c7_c2ab] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond <= VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond;
     t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue;
     t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output := t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2256_c7_e6a8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2256_c7_e6a8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2256_c7_e6a8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2256_c7_e6a8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond <= VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond;
     n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue;
     n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output := n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2256_c7_e6a8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- Submodule level 2
     VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_left := VAR_BIN_OP_SR_uxn_opcodes_h_l2259_c11_1037_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;
     -- t8_MUX[uxn_opcodes_h_l2249_c7_1432] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2249_c7_1432_cond <= VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_cond;
     t8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue;
     t8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output := t8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;

     -- n8_MUX[uxn_opcodes_h_l2252_c7_c2ab] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond <= VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond;
     n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue;
     n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output := n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;

     -- BIN_OP_SL[uxn_opcodes_h_l2259_c11_4f50] LATENCY=0
     -- Inputs
     BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_left <= VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_left;
     BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_right <= VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_right;
     -- Outputs
     VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_return_output := BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2252_c7_c2ab] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2252_c7_c2ab] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2252_c7_c2ab] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2252_c7_c2ab] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;

     -- Submodule level 3
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue := VAR_BIN_OP_SL_uxn_opcodes_h_l2259_c11_4f50_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;
     -- t8_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2256_c7_e6a8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output := result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;

     -- n8_MUX[uxn_opcodes_h_l2249_c7_1432] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2249_c7_1432_cond <= VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_cond;
     n8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue;
     n8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output := n8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2249_c7_1432] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2256_c7_e6a8] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_cond;
     tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output := tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2249_c7_1432] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2249_c7_1432] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2249_c7_1432] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2256_c7_e6a8_return_output;
     -- tmp8_MUX[uxn_opcodes_h_l2252_c7_c2ab] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond;
     tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output := tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2252_c7_c2ab] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output := result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- n8_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2252_c7_c2ab_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2249_c7_1432] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_return_output := result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2249_c7_1432] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_cond;
     tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output := tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;

     -- Submodule level 6
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;
     VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse := VAR_tmp8_MUX_uxn_opcodes_h_l2249_c7_1432_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- tmp8_MUX[uxn_opcodes_h_l2236_c2_5e7c] LATENCY=0
     -- Inputs
     tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond <= VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_cond;
     tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue <= VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iftrue;
     tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse <= VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_iffalse;
     -- Outputs
     VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output := tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;

     -- Submodule level 7
     REG_VAR_tmp8 := VAR_tmp8_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2232_l2266_DUPLICATE_340f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2232_l2266_DUPLICATE_340f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_e848(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2236_c2_5e7c_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2232_l2266_DUPLICATE_340f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_e848_uxn_opcodes_h_l2232_l2266_DUPLICATE_340f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_tmp8 <= REG_VAR_tmp8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     tmp8 <= REG_COMB_tmp8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
