-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 38
entity sub_0CLK_64d180f1 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end sub_0CLK_64d180f1;
architecture arch of sub_0CLK_64d180f1 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2479_c6_7b76]
signal BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2479_c2_f647]
signal t8_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l2479_c2_f647]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2479_c2_f647]
signal n8_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2492_c11_c7a5]
signal BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2492_c7_2cbb]
signal t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2492_c7_2cbb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2492_c7_2cbb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2492_c7_2cbb]
signal result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2492_c7_2cbb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2492_c7_2cbb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2492_c7_2cbb]
signal n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2495_c11_b330]
signal BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l2495_c7_5a92]
signal t8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2495_c7_5a92]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2495_c7_5a92]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2495_c7_5a92]
signal result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2495_c7_5a92]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2495_c7_5a92]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2495_c7_5a92]
signal n8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2498_c11_60ee]
signal BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2498_c7_733d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2498_c7_733d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2498_c7_733d]
signal result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2498_c7_733d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2498_c7_733d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l2498_c7_733d]
signal n8_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2500_c30_b9be]
signal sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_return_output : signed(3 downto 0);

-- BIN_OP_MINUS[uxn_opcodes_h_l2503_c21_3b90]
signal BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_left : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_right : unsigned(7 downto 0);
signal BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_c580( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : signed;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_opc_done := ref_toks_1;
      base.is_vram_write := ref_toks_2;
      base.is_ram_write := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.u8_value := ref_toks_6;
      base.sp_relative_shift := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_pc_updated := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76
BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_left,
BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_right,
BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output);

-- t8_MUX_uxn_opcodes_h_l2479_c2_f647
t8_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
t8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
t8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
t8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647
result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647
result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647
result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647
result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647
result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647
result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647
result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- n8_MUX_uxn_opcodes_h_l2479_c2_f647
n8_MUX_uxn_opcodes_h_l2479_c2_f647 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2479_c2_f647_cond,
n8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue,
n8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse,
n8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5
BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_left,
BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_right,
BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output);

-- t8_MUX_uxn_opcodes_h_l2492_c7_2cbb
t8_MUX_uxn_opcodes_h_l2492_c7_2cbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond,
t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue,
t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse,
t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb
result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb
result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond,
result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb
result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb
result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output);

-- n8_MUX_uxn_opcodes_h_l2492_c7_2cbb
n8_MUX_uxn_opcodes_h_l2492_c7_2cbb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond,
n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue,
n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse,
n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330
BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_left,
BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_right,
BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output);

-- t8_MUX_uxn_opcodes_h_l2495_c7_5a92
t8_MUX_uxn_opcodes_h_l2495_c7_5a92 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond,
t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue,
t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse,
t8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92
result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_cond,
result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92
result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output);

-- n8_MUX_uxn_opcodes_h_l2495_c7_5a92
n8_MUX_uxn_opcodes_h_l2495_c7_5a92 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond,
n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue,
n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse,
n8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee
BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_left,
BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_right,
BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d
result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d
result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_cond,
result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d
result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d
result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_return_output);

-- n8_MUX_uxn_opcodes_h_l2498_c7_733d
n8_MUX_uxn_opcodes_h_l2498_c7_733d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2498_c7_733d_cond,
n8_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue,
n8_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse,
n8_MUX_uxn_opcodes_h_l2498_c7_733d_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be
sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_ins,
sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_x,
sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_y,
sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_return_output);

-- BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90
BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90 : entity work.BIN_OP_MINUS_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_left,
BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_right,
BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output,
 t8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 n8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output,
 t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output,
 n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output,
 t8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output,
 n8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_return_output,
 n8_MUX_uxn_opcodes_h_l2498_c7_733d_return_output,
 sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_return_output,
 BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2489_c3_4109 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l2484_c3_5eed : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2493_c3_d371 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2502_c3_fca8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2495_l2479_l2498_l2492_DUPLICATE_cbdb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_495b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_855d_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_4bb7_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2495_l2498_DUPLICATE_9f3e_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2507_l2475_DUPLICATE_5fde_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2493_c3_d371 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2493_c3_d371;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2502_c3_fca8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2502_c3_fca8;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_right := to_unsigned(2, 2);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue := to_unsigned(1, 1);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2489_c3_4109 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2489_c3_4109;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue := to_unsigned(1, 1);
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_y := resize(to_signed(-1, 2), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l2484_c3_5eed := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l2484_c3_5eed;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_right := to_unsigned(3, 2);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_left := VAR_phase;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse := t8;
     -- BIN_OP_MINUS[uxn_opcodes_h_l2503_c21_3b90] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_left <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_left;
     BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_right <= VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_return_output := BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2495_c11_b330] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_left;
     BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output := BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2498_c11_60ee] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_left;
     BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output := BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_4bb7 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_4bb7_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2492_c11_c7a5] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_left;
     BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output := BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_855d LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_855d_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l2479_c6_7b76] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_left;
     BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output := BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2500_c30_b9be] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_ins;
     sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_x;
     sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_return_output := sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2479_c2_f647_return_output := result.is_ram_write;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2479_c2_f647_return_output := result.is_vram_write;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_495b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_495b_return_output := result.is_opc_done;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2479_c2_f647_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2495_l2479_l2498_l2492_DUPLICATE_cbdb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2495_l2479_l2498_l2492_DUPLICATE_cbdb_return_output := result.u8_value;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2479_c2_f647_return_output := result.is_pc_updated;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2495_l2498_DUPLICATE_9f3e LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2495_l2498_DUPLICATE_9f3e_return_output := result.stack_address_sp_offset;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2479_c6_7b76_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2492_c11_c7a5_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2495_c11_b330_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2498_c11_60ee_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue := VAR_BIN_OP_MINUS_uxn_opcodes_h_l2503_c21_3b90_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_4bb7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_4bb7_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_4bb7_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_495b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_495b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_495b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_855d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_855d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2495_l2498_l2492_DUPLICATE_855d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2495_l2498_DUPLICATE_9f3e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2495_l2498_DUPLICATE_9f3e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2495_l2479_l2498_l2492_DUPLICATE_cbdb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2495_l2479_l2498_l2492_DUPLICATE_cbdb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2495_l2479_l2498_l2492_DUPLICATE_cbdb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2495_l2479_l2498_l2492_DUPLICATE_cbdb_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l2479_c2_f647_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l2479_c2_f647_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l2479_c2_f647_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l2479_c2_f647_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2500_c30_b9be_return_output;
     -- t8_MUX[uxn_opcodes_h_l2495_c7_5a92] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond <= VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond;
     t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue;
     t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output := t8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2498_c7_733d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2498_c7_733d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_return_output := result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2498_c7_733d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2498_c7_733d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;

     -- n8_MUX[uxn_opcodes_h_l2498_c7_733d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2498_c7_733d_cond <= VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_cond;
     n8_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue;
     n8_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_return_output := n8_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2498_c7_733d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;

     -- Submodule level 2
     VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2498_c7_733d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;
     -- t8_MUX[uxn_opcodes_h_l2492_c7_2cbb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond <= VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond;
     t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue;
     t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output := t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2495_c7_5a92] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2495_c7_5a92] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2495_c7_5a92] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2495_c7_5a92] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output := result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2495_c7_5a92] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;

     -- n8_MUX[uxn_opcodes_h_l2495_c7_5a92] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond <= VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_cond;
     n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iftrue;
     n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output := n8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2495_c7_5a92_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2492_c7_2cbb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;

     -- t8_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     t8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     t8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := t8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2492_c7_2cbb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2492_c7_2cbb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output := result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2492_c7_2cbb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;

     -- n8_MUX[uxn_opcodes_h_l2492_c7_2cbb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond <= VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond;
     n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue;
     n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output := n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2492_c7_2cbb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2492_c7_2cbb_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- n8_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     n8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     n8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := n8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2479_c2_f647] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2479_c2_f647_return_output;
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2507_l2475_DUPLICATE_5fde LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2507_l2475_DUPLICATE_5fde_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_c580(
     result,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l2479_c2_f647_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l2479_c2_f647_return_output);

     -- Submodule level 6
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2507_l2475_DUPLICATE_5fde_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_c580_uxn_opcodes_h_l2507_l2475_DUPLICATE_5fde_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
