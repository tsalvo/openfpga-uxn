-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 44
entity and_0CLK_bacf6a1d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end and_0CLK_bacf6a1d;
architecture arch of and_0CLK_bacf6a1d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l877_c6_cb52]
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l877_c1_6daf]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l877_c2_15a8]
signal t8_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l877_c2_15a8]
signal n8_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l877_c2_15a8]
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c2_15a8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l877_c2_15a8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l877_c2_15a8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l877_c2_15a8]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l877_c2_15a8]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l878_c3_6c54[uxn_opcodes_h_l878_c3_6c54]
signal printf_uxn_opcodes_h_l878_c3_6c54_uxn_opcodes_h_l878_c3_6c54_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l882_c11_cd92]
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l882_c7_625f]
signal t8_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l882_c7_625f]
signal n8_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l882_c7_625f]
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l882_c7_625f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l882_c7_625f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l882_c7_625f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l882_c7_625f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l882_c7_625f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l885_c11_2c3d]
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l885_c7_d244]
signal t8_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l885_c7_d244]
signal n8_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l885_c7_d244]
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l885_c7_d244]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l885_c7_d244]
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l885_c7_d244]
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l885_c7_d244]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l885_c7_d244]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l888_c11_3bfa]
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l888_c7_508e]
signal n8_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l888_c7_508e]
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l888_c7_508e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l888_c7_508e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l888_c7_508e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l888_c7_508e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l888_c7_508e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l891_c30_0d52]
signal sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_return_output : signed(3 downto 0);

-- BIN_OP_AND[uxn_opcodes_h_l894_c21_8bfe]
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_left : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_right : unsigned(7 downto 0);
signal BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l896_c11_22ee]
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l896_c7_44a2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l896_c7_44a2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l896_c7_44a2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52
BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_left,
BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_right,
BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_return_output);

-- t8_MUX_uxn_opcodes_h_l877_c2_15a8
t8_MUX_uxn_opcodes_h_l877_c2_15a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l877_c2_15a8_cond,
t8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue,
t8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse,
t8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

-- n8_MUX_uxn_opcodes_h_l877_c2_15a8
n8_MUX_uxn_opcodes_h_l877_c2_15a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l877_c2_15a8_cond,
n8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue,
n8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse,
n8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8
result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_cond,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

-- printf_uxn_opcodes_h_l878_c3_6c54_uxn_opcodes_h_l878_c3_6c54
printf_uxn_opcodes_h_l878_c3_6c54_uxn_opcodes_h_l878_c3_6c54 : entity work.printf_uxn_opcodes_h_l878_c3_6c54_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l878_c3_6c54_uxn_opcodes_h_l878_c3_6c54_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92
BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_left,
BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_right,
BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output);

-- t8_MUX_uxn_opcodes_h_l882_c7_625f
t8_MUX_uxn_opcodes_h_l882_c7_625f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l882_c7_625f_cond,
t8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue,
t8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse,
t8_MUX_uxn_opcodes_h_l882_c7_625f_return_output);

-- n8_MUX_uxn_opcodes_h_l882_c7_625f
n8_MUX_uxn_opcodes_h_l882_c7_625f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l882_c7_625f_cond,
n8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue,
n8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse,
n8_MUX_uxn_opcodes_h_l882_c7_625f_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f
result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_cond,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d
BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_left,
BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_right,
BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output);

-- t8_MUX_uxn_opcodes_h_l885_c7_d244
t8_MUX_uxn_opcodes_h_l885_c7_d244 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l885_c7_d244_cond,
t8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue,
t8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse,
t8_MUX_uxn_opcodes_h_l885_c7_d244_return_output);

-- n8_MUX_uxn_opcodes_h_l885_c7_d244
n8_MUX_uxn_opcodes_h_l885_c7_d244 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l885_c7_d244_cond,
n8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue,
n8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse,
n8_MUX_uxn_opcodes_h_l885_c7_d244_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244
result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_cond,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa
BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_left,
BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_right,
BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output);

-- n8_MUX_uxn_opcodes_h_l888_c7_508e
n8_MUX_uxn_opcodes_h_l888_c7_508e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l888_c7_508e_cond,
n8_MUX_uxn_opcodes_h_l888_c7_508e_iftrue,
n8_MUX_uxn_opcodes_h_l888_c7_508e_iffalse,
n8_MUX_uxn_opcodes_h_l888_c7_508e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e
result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_cond,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output);

-- sp_relative_shift_uxn_opcodes_h_l891_c30_0d52
sp_relative_shift_uxn_opcodes_h_l891_c30_0d52 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_ins,
sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_x,
sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_y,
sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_return_output);

-- BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe
BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe : entity work.BIN_OP_AND_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_left,
BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_right,
BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee
BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_left,
BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_right,
BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_return_output,
 t8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
 n8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output,
 t8_MUX_uxn_opcodes_h_l882_c7_625f_return_output,
 n8_MUX_uxn_opcodes_h_l882_c7_625f_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output,
 t8_MUX_uxn_opcodes_h_l885_c7_d244_return_output,
 n8_MUX_uxn_opcodes_h_l885_c7_d244_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output,
 n8_MUX_uxn_opcodes_h_l888_c7_508e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output,
 sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_return_output,
 BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_679c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l878_c3_6c54_uxn_opcodes_h_l878_c3_6c54_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_397c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_6b8c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_d034_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_6fd2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_3329_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_b60c_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l882_l896_l885_l888_DUPLICATE_75cb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_e84e_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l902_l873_DUPLICATE_17ae_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_right := to_unsigned(4, 3);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_6b8c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l893_c3_6b8c;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_y := resize(to_signed(-1, 2), 4);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iffalse := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_397c := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l883_c3_397c;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_679c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l879_c3_679c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_right := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_left := VAR_phase;
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l888_c11_3bfa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_left;
     BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output := BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_b60c LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_b60c_return_output := result.sp_relative_shift;

     -- BIN_OP_AND[uxn_opcodes_h_l894_c21_8bfe] LATENCY=0
     -- Inputs
     BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_left <= VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_left;
     BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_right <= VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_right;
     -- Outputs
     VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_return_output := BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l882_l896_l885_l888_DUPLICATE_75cb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l882_l896_l885_l888_DUPLICATE_75cb_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l877_c6_cb52] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_left;
     BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output := BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_3329 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_3329_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l882_c11_cd92] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_left;
     BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output := BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l885_c11_2c3d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_left;
     BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output := BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_e84e LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_e84e_return_output := result.stack_address_sp_offset;

     -- sp_relative_shift[uxn_opcodes_h_l891_c30_0d52] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_ins;
     sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_x <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_x;
     sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_y <= VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_return_output := sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_6fd2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_6fd2_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l896_c11_22ee] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_left;
     BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output := BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_d034 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_d034_return_output := result.u8_value;

     -- Submodule level 1
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iftrue := VAR_BIN_OP_AND_uxn_opcodes_h_l894_c21_8bfe_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l877_c6_cb52_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l882_c11_cd92_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l885_c11_2c3d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l888_c11_3bfa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l896_c11_22ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_b60c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_b60c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_b60c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_b60c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l882_l896_l885_l888_DUPLICATE_75cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l882_l896_l885_l888_DUPLICATE_75cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l882_l896_l885_l888_DUPLICATE_75cb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l882_l896_l885_l888_DUPLICATE_75cb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_6fd2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_6fd2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_6fd2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_6fd2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_3329_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_3329_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_3329_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l882_l896_l885_l877_DUPLICATE_3329_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_e84e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l885_l888_DUPLICATE_e84e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_d034_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_d034_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_d034_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l882_l885_l877_l888_DUPLICATE_d034_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l891_c30_0d52_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l896_c7_44a2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_return_output;

     -- t8_MUX[uxn_opcodes_h_l885_c7_d244] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l885_c7_d244_cond <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_cond;
     t8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue;
     t8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_return_output := t8_MUX_uxn_opcodes_h_l885_c7_d244_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l877_c1_6daf] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l896_c7_44a2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l888_c7_508e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_return_output := result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_return_output;

     -- n8_MUX[uxn_opcodes_h_l888_c7_508e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l888_c7_508e_cond <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_cond;
     n8_MUX_uxn_opcodes_h_l888_c7_508e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_iftrue;
     n8_MUX_uxn_opcodes_h_l888_c7_508e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_return_output := n8_MUX_uxn_opcodes_h_l888_c7_508e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l896_c7_44a2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l888_c7_508e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l888_c7_508e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_return_output;

     -- Submodule level 2
     VAR_printf_uxn_opcodes_h_l878_c3_6c54_uxn_opcodes_h_l878_c3_6c54_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l877_c1_6daf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse := VAR_n8_MUX_uxn_opcodes_h_l888_c7_508e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l896_c7_44a2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l896_c7_44a2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l896_c7_44a2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l888_c7_508e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l888_c7_508e_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse := VAR_t8_MUX_uxn_opcodes_h_l885_c7_d244_return_output;
     -- n8_MUX[uxn_opcodes_h_l885_c7_d244] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l885_c7_d244_cond <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_cond;
     n8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_iftrue;
     n8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_return_output := n8_MUX_uxn_opcodes_h_l885_c7_d244_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l885_c7_d244] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l885_c7_d244] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l888_c7_508e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l888_c7_508e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_return_output;

     -- t8_MUX[uxn_opcodes_h_l882_c7_625f] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l882_c7_625f_cond <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_cond;
     t8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue;
     t8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_return_output := t8_MUX_uxn_opcodes_h_l882_c7_625f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l888_c7_508e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l885_c7_d244] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_cond;
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_return_output := result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_return_output;

     -- printf_uxn_opcodes_h_l878_c3_6c54[uxn_opcodes_h_l878_c3_6c54] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l878_c3_6c54_uxn_opcodes_h_l878_c3_6c54_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l878_c3_6c54_uxn_opcodes_h_l878_c3_6c54_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse := VAR_n8_MUX_uxn_opcodes_h_l885_c7_d244_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l888_c7_508e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l888_c7_508e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l888_c7_508e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l885_c7_d244_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l885_c7_d244_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse := VAR_t8_MUX_uxn_opcodes_h_l882_c7_625f_return_output;
     -- n8_MUX[uxn_opcodes_h_l882_c7_625f] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l882_c7_625f_cond <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_cond;
     n8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_iftrue;
     n8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_return_output := n8_MUX_uxn_opcodes_h_l882_c7_625f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l882_c7_625f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l885_c7_d244] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l885_c7_d244] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l882_c7_625f] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_cond;
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_return_output := result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l885_c7_d244] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l882_c7_625f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output;

     -- t8_MUX[uxn_opcodes_h_l877_c2_15a8] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l877_c2_15a8_cond <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_cond;
     t8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue;
     t8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output := t8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse := VAR_n8_MUX_uxn_opcodes_h_l882_c7_625f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l885_c7_d244_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l885_c7_d244_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l885_c7_d244_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l882_c7_625f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l882_c7_625f_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l877_c2_15a8] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;

     -- n8_MUX[uxn_opcodes_h_l877_c2_15a8] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l877_c2_15a8_cond <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_cond;
     n8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue;
     n8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output := n8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l882_c7_625f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l882_c7_625f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l877_c2_15a8] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_cond;
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_return_output := result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l877_c2_15a8] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l882_c7_625f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l882_c7_625f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l882_c7_625f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l882_c7_625f_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l877_c2_15a8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l877_c2_15a8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l877_c2_15a8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l902_l873_DUPLICATE_17ae LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l902_l873_DUPLICATE_17ae_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l877_c2_15a8_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l877_c2_15a8_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l902_l873_DUPLICATE_17ae_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l902_l873_DUPLICATE_17ae_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
