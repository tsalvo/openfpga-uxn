-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 53
entity gth_0CLK_6d7675a8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_6d7675a8;
architecture arch of gth_0CLK_6d7675a8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1921_c6_260b]
signal BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1921_c1_0118]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1921_c2_5b9d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1921_c2_5b9d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1921_c2_5b9d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1921_c2_5b9d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1921_c2_5b9d]
signal result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1921_c2_5b9d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1921_c2_5b9d]
signal t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1921_c2_5b9d]
signal n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1922_c3_f007[uxn_opcodes_h_l1922_c3_f007]
signal printf_uxn_opcodes_h_l1922_c3_f007_uxn_opcodes_h_l1922_c3_f007_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1926_c11_843f]
signal BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1926_c7_e2c4]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1926_c7_e2c4]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1926_c7_e2c4]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1926_c7_e2c4]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1926_c7_e2c4]
signal result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1926_c7_e2c4]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1926_c7_e2c4]
signal t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1926_c7_e2c4]
signal n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1929_c11_ba82]
signal BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1929_c7_327d]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1929_c7_327d]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1929_c7_327d]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1929_c7_327d]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1929_c7_327d]
signal result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1929_c7_327d]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1929_c7_327d]
signal t8_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1929_c7_327d]
signal n8_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1933_c11_c594]
signal BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1933_c7_a849]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1933_c7_a849]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1933_c7_a849]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1933_c7_a849]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1933_c7_a849]
signal result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1933_c7_a849]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1933_c7_a849]
signal n8_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1936_c11_738a]
signal BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1936_c7_fdb2]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1936_c7_fdb2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1936_c7_fdb2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1936_c7_fdb2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1936_c7_fdb2]
signal result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(7 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1936_c7_fdb2]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : signed(3 downto 0);

-- n8_MUX[uxn_opcodes_h_l1936_c7_fdb2]
signal n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1939_c30_5867]
signal sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1942_c21_5b3e]
signal BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1942_c21_81f7]
signal MUX_uxn_opcodes_h_l1942_c21_81f7_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1942_c21_81f7_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1942_c21_81f7_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1942_c21_81f7_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1944_c11_cb7a]
signal BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1944_c7_d9d8]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1944_c7_d9d8]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1944_c7_d9d8]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_641b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.u8_value := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b
BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_left,
BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_right,
BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d
result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

-- t8_MUX_uxn_opcodes_h_l1921_c2_5b9d
t8_MUX_uxn_opcodes_h_l1921_c2_5b9d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond,
t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue,
t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse,
t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

-- n8_MUX_uxn_opcodes_h_l1921_c2_5b9d
n8_MUX_uxn_opcodes_h_l1921_c2_5b9d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond,
n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue,
n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse,
n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

-- printf_uxn_opcodes_h_l1922_c3_f007_uxn_opcodes_h_l1922_c3_f007
printf_uxn_opcodes_h_l1922_c3_f007_uxn_opcodes_h_l1922_c3_f007 : entity work.printf_uxn_opcodes_h_l1922_c3_f007_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1922_c3_f007_uxn_opcodes_h_l1922_c3_f007_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f
BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_left,
BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_right,
BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4
result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4
result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4
result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4
result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond,
result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4
result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output);

-- t8_MUX_uxn_opcodes_h_l1926_c7_e2c4
t8_MUX_uxn_opcodes_h_l1926_c7_e2c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond,
t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue,
t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse,
t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output);

-- n8_MUX_uxn_opcodes_h_l1926_c7_e2c4
n8_MUX_uxn_opcodes_h_l1926_c7_e2c4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond,
n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue,
n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse,
n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82
BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_left,
BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_right,
BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d
result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d
result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d
result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d
result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_cond,
result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d
result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output);

-- t8_MUX_uxn_opcodes_h_l1929_c7_327d
t8_MUX_uxn_opcodes_h_l1929_c7_327d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1929_c7_327d_cond,
t8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue,
t8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse,
t8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output);

-- n8_MUX_uxn_opcodes_h_l1929_c7_327d
n8_MUX_uxn_opcodes_h_l1929_c7_327d : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1929_c7_327d_cond,
n8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue,
n8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse,
n8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594
BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_left,
BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_right,
BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849
result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849
result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849
result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849
result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_cond,
result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849
result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output);

-- n8_MUX_uxn_opcodes_h_l1933_c7_a849
n8_MUX_uxn_opcodes_h_l1933_c7_a849 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1933_c7_a849_cond,
n8_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue,
n8_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse,
n8_MUX_uxn_opcodes_h_l1933_c7_a849_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a
BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_left,
BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_right,
BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2
result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2
result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2
result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2
result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond,
result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2
result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output);

-- n8_MUX_uxn_opcodes_h_l1936_c7_fdb2
n8_MUX_uxn_opcodes_h_l1936_c7_fdb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond,
n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue,
n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse,
n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1939_c30_5867
sp_relative_shift_uxn_opcodes_h_l1939_c30_5867 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_ins,
sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_x,
sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_y,
sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e
BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_left,
BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_right,
BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_return_output);

-- MUX_uxn_opcodes_h_l1942_c21_81f7
MUX_uxn_opcodes_h_l1942_c21_81f7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1942_c21_81f7_cond,
MUX_uxn_opcodes_h_l1942_c21_81f7_iftrue,
MUX_uxn_opcodes_h_l1942_c21_81f7_iffalse,
MUX_uxn_opcodes_h_l1942_c21_81f7_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a
BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_left,
BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_right,
BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8
result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8
result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8
result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
 t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
 n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output,
 t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output,
 n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output,
 t8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output,
 n8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output,
 n8_MUX_uxn_opcodes_h_l1933_c7_a849_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output,
 n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output,
 sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_return_output,
 MUX_uxn_opcodes_h_l1942_c21_81f7_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iffalse : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1923_c3_395b : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1922_c3_f007_uxn_opcodes_h_l1922_c3_f007_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1927_c3_183c : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1931_c3_2333 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1934_c3_4db9 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1941_c3_1759 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1936_c7_fdb2_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_a41b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_cb9c_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_104a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_37d9_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1926_l1944_l1936_l1933_l1929_DUPLICATE_b74b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1917_l1950_DUPLICATE_e86e_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1941_c3_1759 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1941_c3_1759;
     VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_right := to_unsigned(2, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1931_c3_2333 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1931_c3_2333;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1927_c3_183c := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1927_c3_183c;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_right := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1923_c3_395b := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1923_c3_395b;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1934_c3_4db9 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1934_c3_4db9;
     VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_right := to_unsigned(3, 2);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iffalse := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1926_l1944_l1936_l1933_l1929_DUPLICATE_b74b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1926_l1944_l1936_l1933_l1929_DUPLICATE_b74b_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l1936_c11_738a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_a41b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_a41b_return_output := result.is_sp_shift;

     -- BIN_OP_GT[uxn_opcodes_h_l1942_c21_5b3e] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_left;
     BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_return_output := BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_37d9 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_37d9_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1926_c11_843f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1944_c11_cb7a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1929_c11_ba82] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_left;
     BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output := BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1939_c30_5867] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_ins;
     sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_x;
     sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_return_output := sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_104a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_104a_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1921_c6_260b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_left;
     BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output := BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_cb9c LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_cb9c_return_output := result.is_stack_write;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l1936_c7_fdb2] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1936_c7_fdb2_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1933_c11_c594] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_left;
     BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output := BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1921_c6_260b_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1926_c11_843f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1929_c11_ba82_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1933_c11_c594_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1936_c11_738a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1944_c11_cb7a_return_output;
     VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1942_c21_5b3e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_37d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_37d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_37d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_37d9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_37d9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1926_l1944_l1936_l1933_l1929_DUPLICATE_b74b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1926_l1944_l1936_l1933_l1929_DUPLICATE_b74b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1926_l1944_l1936_l1933_l1929_DUPLICATE_b74b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1926_l1944_l1936_l1933_l1929_DUPLICATE_b74b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1926_l1944_l1936_l1933_l1929_DUPLICATE_b74b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_a41b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_a41b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_a41b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_a41b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_a41b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_cb9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_cb9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_cb9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_cb9c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1926_l1921_l1944_l1933_l1929_DUPLICATE_cb9c_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_104a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_104a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_104a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_104a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1926_l1921_l1936_l1933_l1929_DUPLICATE_104a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1936_c7_fdb2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1939_c30_5867_return_output;
     -- MUX[uxn_opcodes_h_l1942_c21_81f7] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1942_c21_81f7_cond <= VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_cond;
     MUX_uxn_opcodes_h_l1942_c21_81f7_iftrue <= VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_iftrue;
     MUX_uxn_opcodes_h_l1942_c21_81f7_iffalse <= VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_return_output := MUX_uxn_opcodes_h_l1942_c21_81f7_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1944_c7_d9d8] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output;

     -- n8_MUX[uxn_opcodes_h_l1936_c7_fdb2] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond <= VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond;
     n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue;
     n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output := n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1944_c7_d9d8] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output;

     -- t8_MUX[uxn_opcodes_h_l1929_c7_327d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1929_c7_327d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_cond;
     t8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue;
     t8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output := t8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1921_c1_0118] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1944_c7_d9d8] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1936_c7_fdb2] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1936_c7_fdb2] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue := VAR_MUX_uxn_opcodes_h_l1942_c21_81f7_return_output;
     VAR_printf_uxn_opcodes_h_l1922_c3_f007_uxn_opcodes_h_l1922_c3_f007_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1921_c1_0118_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1944_c7_d9d8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1936_c7_fdb2] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output := result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;

     -- n8_MUX[uxn_opcodes_h_l1933_c7_a849] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1933_c7_a849_cond <= VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_cond;
     n8_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue;
     n8_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_return_output := n8_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1936_c7_fdb2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1933_c7_a849] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1936_c7_fdb2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;

     -- t8_MUX[uxn_opcodes_h_l1926_c7_e2c4] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond <= VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond;
     t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue;
     t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output := t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;

     -- printf_uxn_opcodes_h_l1922_c3_f007[uxn_opcodes_h_l1922_c3_f007] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1922_c3_f007_uxn_opcodes_h_l1922_c3_f007_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1922_c3_f007_uxn_opcodes_h_l1922_c3_f007_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1933_c7_a849] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1936_c7_fdb2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1936_c7_fdb2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1929_c7_327d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1933_c7_a849] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1929_c7_327d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1933_c7_a849] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1933_c7_a849] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;

     -- n8_MUX[uxn_opcodes_h_l1929_c7_327d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1929_c7_327d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_cond;
     n8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue;
     n8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output := n8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1933_c7_a849] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_return_output := result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;

     -- t8_MUX[uxn_opcodes_h_l1921_c2_5b9d] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond <= VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond;
     t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue;
     t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output := t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1933_c7_a849_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;
     -- n8_MUX[uxn_opcodes_h_l1926_c7_e2c4] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond <= VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond;
     n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue;
     n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output := n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1929_c7_327d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1929_c7_327d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1929_c7_327d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1926_c7_e2c4] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1926_c7_e2c4] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1929_c7_327d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1929_c7_327d_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1926_c7_e2c4] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1926_c7_e2c4] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output := result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1926_c7_e2c4] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;

     -- n8_MUX[uxn_opcodes_h_l1921_c2_5b9d] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond <= VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond;
     n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue;
     n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output := n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1921_c2_5b9d] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1926_c7_e2c4] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1921_c2_5b9d] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1926_c7_e2c4_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1921_c2_5b9d] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1921_c2_5b9d] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1921_c2_5b9d] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1921_c2_5b9d] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output := result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1917_l1950_DUPLICATE_e86e LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1917_l1950_DUPLICATE_e86e_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_641b(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1921_c2_5b9d_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1917_l1950_DUPLICATE_e86e_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_641b_uxn_opcodes_h_l1917_l1950_DUPLICATE_e86e_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
