-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity equ_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end equ_0CLK_85d5529e;
architecture arch of equ_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1114_c6_fee9]
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1114_c1_db31]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1114_c2_f453]
signal n8_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1114_c2_f453]
signal t8_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1114_c2_f453]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1114_c2_f453]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1114_c2_f453]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1114_c2_f453]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1114_c2_f453]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1114_c2_f453]
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(7 downto 0);

-- printf_uxn_opcodes_h_l1115_c3_d457[uxn_opcodes_h_l1115_c3_d457]
signal printf_uxn_opcodes_h_l1115_c3_d457_uxn_opcodes_h_l1115_c3_d457_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1119_c11_52e0]
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1119_c7_946e]
signal n8_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1119_c7_946e]
signal t8_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1119_c7_946e]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1119_c7_946e]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1119_c7_946e]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1119_c7_946e]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1119_c7_946e]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1119_c7_946e]
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1122_c11_f7b9]
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1122_c7_7af3]
signal n8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l1122_c7_7af3]
signal t8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1122_c7_7af3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1122_c7_7af3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1122_c7_7af3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1122_c7_7af3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1122_c7_7af3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1122_c7_7af3]
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1125_c11_7d28]
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1125_c7_0636]
signal n8_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1125_c7_0636]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1125_c7_0636]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1125_c7_0636]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1125_c7_0636]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1125_c7_0636]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1125_c7_0636]
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(7 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1128_c30_f3d2]
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1131_c21_9764]
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1131_c21_8345]
signal MUX_uxn_opcodes_h_l1131_c21_8345_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_8345_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_8345_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1131_c21_8345_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1133_c11_83ed]
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1133_c7_5192]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1133_c7_5192]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1133_c7_5192]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5b93( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_stack_write := ref_toks_1;
      base.stack_address_sp_offset := ref_toks_2;
      base.is_sp_shift := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.u8_value := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_left,
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_right,
BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_return_output);

-- n8_MUX_uxn_opcodes_h_l1114_c2_f453
n8_MUX_uxn_opcodes_h_l1114_c2_f453 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1114_c2_f453_cond,
n8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue,
n8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse,
n8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

-- t8_MUX_uxn_opcodes_h_l1114_c2_f453
t8_MUX_uxn_opcodes_h_l1114_c2_f453 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1114_c2_f453_cond,
t8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue,
t8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse,
t8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_cond,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

-- printf_uxn_opcodes_h_l1115_c3_d457_uxn_opcodes_h_l1115_c3_d457
printf_uxn_opcodes_h_l1115_c3_d457_uxn_opcodes_h_l1115_c3_d457 : entity work.printf_uxn_opcodes_h_l1115_c3_d457_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1115_c3_d457_uxn_opcodes_h_l1115_c3_d457_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_left,
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_right,
BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output);

-- n8_MUX_uxn_opcodes_h_l1119_c7_946e
n8_MUX_uxn_opcodes_h_l1119_c7_946e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1119_c7_946e_cond,
n8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue,
n8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse,
n8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output);

-- t8_MUX_uxn_opcodes_h_l1119_c7_946e
t8_MUX_uxn_opcodes_h_l1119_c7_946e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1119_c7_946e_cond,
t8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue,
t8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse,
t8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_cond,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_left,
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_right,
BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output);

-- n8_MUX_uxn_opcodes_h_l1122_c7_7af3
n8_MUX_uxn_opcodes_h_l1122_c7_7af3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond,
n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue,
n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse,
n8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output);

-- t8_MUX_uxn_opcodes_h_l1122_c7_7af3
t8_MUX_uxn_opcodes_h_l1122_c7_7af3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond,
t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue,
t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse,
t8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_left,
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_right,
BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output);

-- n8_MUX_uxn_opcodes_h_l1125_c7_0636
n8_MUX_uxn_opcodes_h_l1125_c7_0636 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1125_c7_0636_cond,
n8_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue,
n8_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse,
n8_MUX_uxn_opcodes_h_l1125_c7_0636_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_cond,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2
sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_ins,
sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_x,
sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_y,
sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_left,
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_right,
BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_return_output);

-- MUX_uxn_opcodes_h_l1131_c21_8345
MUX_uxn_opcodes_h_l1131_c21_8345 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1131_c21_8345_cond,
MUX_uxn_opcodes_h_l1131_c21_8345_iftrue,
MUX_uxn_opcodes_h_l1131_c21_8345_iffalse,
MUX_uxn_opcodes_h_l1131_c21_8345_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_left,
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_right,
BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_return_output,
 n8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
 t8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output,
 n8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output,
 t8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output,
 n8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output,
 t8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output,
 n8_MUX_uxn_opcodes_h_l1125_c7_0636_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_return_output,
 sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_return_output,
 MUX_uxn_opcodes_h_l1131_c21_8345_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iffalse : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_055f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1115_c3_d457_uxn_opcodes_h_l1115_c3_d457_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_eaa8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_4b54 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_8345_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_8345_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_8345_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1131_c21_8345_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_93d1_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_cd31_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_45bd_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_0d24_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_fdea_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_239a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1139_l1110_DUPLICATE_5556_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_4b54 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1130_c3_4b54;
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iffalse := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1131_c21_8345_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1131_c21_8345_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue := to_unsigned(1, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_eaa8 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1120_c3_eaa8;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_y := resize(to_signed(-1, 2), 4);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_right := to_unsigned(3, 2);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_055f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1116_c3_055f;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_93d1 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_93d1_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_0d24 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_0d24_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1122_c11_f7b9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1128_c30_f3d2] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_ins;
     sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_x;
     sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_return_output := sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1133_c11_83ed] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_left;
     BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output := BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_cd31 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_cd31_return_output := result.is_sp_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1119_c11_52e0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_left;
     BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output := BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1125_c11_7d28] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_left;
     BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output := BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1131_c21_9764] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_left;
     BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_return_output := BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_239a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_239a_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_45bd LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_45bd_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1114_c6_fee9] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_left;
     BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output := BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_fdea LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_fdea_return_output := result.is_opc_done;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1114_c6_fee9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1119_c11_52e0_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1122_c11_f7b9_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1125_c11_7d28_return_output;
     VAR_MUX_uxn_opcodes_h_l1131_c21_8345_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1131_c21_9764_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1133_c11_83ed_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_45bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_45bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_45bd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_45bd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_fdea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_fdea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_fdea_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1125_l1119_l1133_l1122_DUPLICATE_fdea_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_cd31_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_cd31_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_cd31_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_cd31_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_93d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_93d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_93d1_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1114_l1119_l1133_l1122_DUPLICATE_93d1_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_239a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1125_l1122_DUPLICATE_239a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_0d24_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_0d24_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_0d24_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1114_l1125_l1119_l1122_DUPLICATE_0d24_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1128_c30_f3d2_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1125_c7_0636] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1133_c7_5192] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1133_c7_5192] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_return_output;

     -- n8_MUX[uxn_opcodes_h_l1125_c7_0636] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1125_c7_0636_cond <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_cond;
     n8_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue;
     n8_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_return_output := n8_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1114_c1_db31] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1133_c7_5192] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_return_output;

     -- t8_MUX[uxn_opcodes_h_l1122_c7_7af3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond;
     t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue;
     t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output := t8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;

     -- MUX[uxn_opcodes_h_l1131_c21_8345] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1131_c21_8345_cond <= VAR_MUX_uxn_opcodes_h_l1131_c21_8345_cond;
     MUX_uxn_opcodes_h_l1131_c21_8345_iftrue <= VAR_MUX_uxn_opcodes_h_l1131_c21_8345_iftrue;
     MUX_uxn_opcodes_h_l1131_c21_8345_iffalse <= VAR_MUX_uxn_opcodes_h_l1131_c21_8345_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1131_c21_8345_return_output := MUX_uxn_opcodes_h_l1131_c21_8345_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1125_c7_0636] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue := VAR_MUX_uxn_opcodes_h_l1131_c21_8345_return_output;
     VAR_printf_uxn_opcodes_h_l1115_c3_d457_uxn_opcodes_h_l1115_c3_d457_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1114_c1_db31_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1133_c7_5192_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1133_c7_5192_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1133_c7_5192_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1122_c7_7af3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1125_c7_0636] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1125_c7_0636] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_return_output := result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;

     -- n8_MUX[uxn_opcodes_h_l1122_c7_7af3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_cond;
     n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue;
     n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output := n8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1119_c7_946e] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1119_c7_946e_cond <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_cond;
     t8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue;
     t8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output := t8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1122_c7_7af3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;

     -- printf_uxn_opcodes_h_l1115_c3_d457[uxn_opcodes_h_l1115_c3_d457] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1115_c3_d457_uxn_opcodes_h_l1115_c3_d457_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1115_c3_d457_uxn_opcodes_h_l1115_c3_d457_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1125_c7_0636] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1125_c7_0636] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1125_c7_0636_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1119_c7_946e] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1122_c7_7af3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1122_c7_7af3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1119_c7_946e] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1119_c7_946e_cond <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_cond;
     n8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue;
     n8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output := n8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1122_c7_7af3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1119_c7_946e] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;

     -- t8_MUX[uxn_opcodes_h_l1114_c2_f453] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1114_c2_f453_cond <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_cond;
     t8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue;
     t8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output := t8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1122_c7_7af3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1122_c7_7af3_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1114_c2_f453] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;

     -- n8_MUX[uxn_opcodes_h_l1114_c2_f453] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1114_c2_f453_cond <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_cond;
     n8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue;
     n8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output := n8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1119_c7_946e] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1119_c7_946e] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_return_output := result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1119_c7_946e] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1114_c2_f453] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1119_c7_946e] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1119_c7_946e_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1114_c2_f453] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1114_c2_f453] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1114_c2_f453] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1114_c2_f453] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_return_output := result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1139_l1110_DUPLICATE_5556 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1139_l1110_DUPLICATE_5556_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5b93(
     result,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1114_c2_f453_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1114_c2_f453_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1139_l1110_DUPLICATE_5556_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5b93_uxn_opcodes_h_l1139_l1110_DUPLICATE_5556_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
