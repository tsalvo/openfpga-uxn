-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- -- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 51
entity lth_0CLK_57104a4d is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_57104a4d;
architecture arch of lth_0CLK_57104a4d is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l2007_c6_e274]
signal BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2007_c2_cec3]
signal n8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2007_c2_cec3]
signal t8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2007_c2_cec3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2007_c2_cec3]
signal result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2007_c2_cec3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2007_c2_cec3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2007_c2_cec3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2007_c2_cec3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2012_c11_73e6]
signal BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2012_c7_8196]
signal n8_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2012_c7_8196]
signal t8_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2012_c7_8196]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2012_c7_8196]
signal result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2012_c7_8196]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2012_c7_8196]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2012_c7_8196]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2012_c7_8196]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2015_c11_c0e2]
signal BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2015_c7_e35b]
signal n8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(7 downto 0);

-- t8_MUX[uxn_opcodes_h_l2015_c7_e35b]
signal t8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2015_c7_e35b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2015_c7_e35b]
signal result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2015_c7_e35b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2015_c7_e35b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2015_c7_e35b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2015_c7_e35b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2019_c11_75aa]
signal BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2019_c7_3712]
signal n8_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2019_c7_3712]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2019_c7_3712]
signal result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2019_c7_3712]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2019_c7_3712]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2019_c7_3712]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2019_c7_3712]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2022_c11_25fa]
signal BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l2022_c7_0bd0]
signal n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2022_c7_0bd0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l2022_c7_0bd0]
signal result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2022_c7_0bd0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2022_c7_0bd0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l2022_c7_0bd0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : signed(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2022_c7_0bd0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l2025_c30_37d8]
signal sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l2028_c21_c95b]
signal BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l2028_c21_d191]
signal MUX_uxn_opcodes_h_l2028_c21_d191_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l2028_c21_d191_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2028_c21_d191_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l2028_c21_d191_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l2030_c11_576c]
signal BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l2030_c7_005a]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l2030_c7_005a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l2030_c7_005a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_3345( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed;
 ref_toks_6 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.stack_address_sp_offset := ref_toks_1;
      base.u8_value := ref_toks_2;
      base.is_stack_write := ref_toks_3;
      base.is_opc_done := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;
      base.is_sp_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274
BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_left,
BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_right,
BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output);

-- n8_MUX_uxn_opcodes_h_l2007_c2_cec3
n8_MUX_uxn_opcodes_h_l2007_c2_cec3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond,
n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue,
n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse,
n8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

-- t8_MUX_uxn_opcodes_h_l2007_c2_cec3
t8_MUX_uxn_opcodes_h_l2007_c2_cec3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond,
t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue,
t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse,
t8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3
result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_cond,
result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3
result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3
result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3
result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3
result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6
BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_left,
BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_right,
BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output);

-- n8_MUX_uxn_opcodes_h_l2012_c7_8196
n8_MUX_uxn_opcodes_h_l2012_c7_8196 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2012_c7_8196_cond,
n8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue,
n8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse,
n8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output);

-- t8_MUX_uxn_opcodes_h_l2012_c7_8196
t8_MUX_uxn_opcodes_h_l2012_c7_8196 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2012_c7_8196_cond,
t8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue,
t8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse,
t8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_cond,
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2
BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_left,
BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_right,
BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output);

-- n8_MUX_uxn_opcodes_h_l2015_c7_e35b
n8_MUX_uxn_opcodes_h_l2015_c7_e35b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond,
n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue,
n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse,
n8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output);

-- t8_MUX_uxn_opcodes_h_l2015_c7_e35b
t8_MUX_uxn_opcodes_h_l2015_c7_e35b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond,
t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue,
t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse,
t8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b
result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_cond,
result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b
result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b
result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b
result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b
result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa
BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_left,
BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_right,
BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output);

-- n8_MUX_uxn_opcodes_h_l2019_c7_3712
n8_MUX_uxn_opcodes_h_l2019_c7_3712 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2019_c7_3712_cond,
n8_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue,
n8_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse,
n8_MUX_uxn_opcodes_h_l2019_c7_3712_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_cond,
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa
BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_left,
BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_right,
BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output);

-- n8_MUX_uxn_opcodes_h_l2022_c7_0bd0
n8_MUX_uxn_opcodes_h_l2022_c7_0bd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond,
n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue,
n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse,
n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0
result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond,
result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0
result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0
result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0
result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0
result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output);

-- sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8
sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_ins,
sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_x,
sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_y,
sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b
BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_left,
BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_right,
BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_return_output);

-- MUX_uxn_opcodes_h_l2028_c21_d191
MUX_uxn_opcodes_h_l2028_c21_d191 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l2028_c21_d191_cond,
MUX_uxn_opcodes_h_l2028_c21_d191_iftrue,
MUX_uxn_opcodes_h_l2028_c21_d191_iffalse,
MUX_uxn_opcodes_h_l2028_c21_d191_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c
BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_left,
BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_right,
BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a
result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output,
 n8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
 t8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output,
 n8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output,
 t8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output,
 n8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output,
 t8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output,
 n8_MUX_uxn_opcodes_h_l2019_c7_3712_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output,
 n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output,
 sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_return_output,
 BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_return_output,
 MUX_uxn_opcodes_h_l2028_c21_d191_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2009_c3_3d3f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2013_c3_14e4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2017_c3_a4f3 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2020_c3_358a : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2027_c3_4f8f : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2022_c7_0bd0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2028_c21_d191_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2028_c21_d191_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2028_c21_d191_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l2028_c21_d191_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_582e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_09dc_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_29e8_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_ad28_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2030_DUPLICATE_0e95_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2036_l2003_DUPLICATE_bab3_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2027_c3_4f8f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2027_c3_4f8f;
     VAR_MUX_uxn_opcodes_h_l2028_c21_d191_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2013_c3_14e4 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2013_c3_14e4;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2009_c3_3d3f := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2009_c3_3d3f;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l2028_c21_d191_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_right := to_unsigned(4, 3);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue := to_unsigned(0, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_right := to_unsigned(3, 2);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_right := to_unsigned(5, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2017_c3_a4f3 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2017_c3_a4f3;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_y := resize(to_signed(-1, 2), 4);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2020_c3_358a := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l2020_c3_358a;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l2012_c11_73e6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_left;
     BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output := BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2030_c11_576c] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_left;
     BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output := BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l2025_c30_37d8] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_ins;
     sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_x <= VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_x;
     sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_y <= VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_return_output := sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2007_c6_e274] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_left;
     BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output := BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_ad28 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_ad28_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2030_DUPLICATE_0e95 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2030_DUPLICATE_0e95_return_output := result.is_opc_done;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_29e8 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_29e8_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l2019_c11_75aa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_left;
     BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output := BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output;

     -- result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d[uxn_opcodes_h_l2022_c7_0bd0] LATENCY=0
     VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2022_c7_0bd0_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_582e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_582e_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l2022_c11_25fa] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_left;
     BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output := BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l2015_c11_c0e2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_left;
     BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output := BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;

     -- BIN_OP_LT[uxn_opcodes_h_l2028_c21_c95b] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_left;
     BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_return_output := BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_09dc LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_09dc_return_output := result.is_stack_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2007_c6_e274_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2012_c11_73e6_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2015_c11_c0e2_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2019_c11_75aa_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2022_c11_25fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l2030_c11_576c_return_output;
     VAR_MUX_uxn_opcodes_h_l2028_c21_d191_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l2028_c21_c95b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_29e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_29e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_29e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_29e8_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_29e8_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2030_DUPLICATE_0e95_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2030_DUPLICATE_0e95_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2030_DUPLICATE_0e95_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2030_DUPLICATE_0e95_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2030_DUPLICATE_0e95_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_ad28_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_ad28_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_ad28_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_ad28_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_ad28_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_09dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_09dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_09dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_09dc_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l2019_l2015_l2012_l2007_l2030_DUPLICATE_09dc_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_582e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_582e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_582e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_582e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l2022_l2019_l2015_l2012_l2007_DUPLICATE_582e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse := VAR_result_stack_address_sp_offset_FALSE_INPUT_MUX_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l2022_c7_0bd0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l2025_c30_37d8_return_output;
     -- MUX[uxn_opcodes_h_l2028_c21_d191] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l2028_c21_d191_cond <= VAR_MUX_uxn_opcodes_h_l2028_c21_d191_cond;
     MUX_uxn_opcodes_h_l2028_c21_d191_iftrue <= VAR_MUX_uxn_opcodes_h_l2028_c21_d191_iftrue;
     MUX_uxn_opcodes_h_l2028_c21_d191_iffalse <= VAR_MUX_uxn_opcodes_h_l2028_c21_d191_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l2028_c21_d191_return_output := MUX_uxn_opcodes_h_l2028_c21_d191_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2030_c7_005a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_return_output;

     -- n8_MUX[uxn_opcodes_h_l2022_c7_0bd0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond <= VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond;
     n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue;
     n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output := n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2030_c7_005a] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2030_c7_005a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2022_c7_0bd0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2022_c7_0bd0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2015_c7_e35b] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond <= VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond;
     t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue;
     t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output := t8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue := VAR_MUX_uxn_opcodes_h_l2028_c21_d191_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2030_c7_005a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2030_c7_005a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2030_c7_005a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2022_c7_0bd0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;

     -- t8_MUX[uxn_opcodes_h_l2012_c7_8196] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2012_c7_8196_cond <= VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_cond;
     t8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue;
     t8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output := t8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2022_c7_0bd0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output := result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2022_c7_0bd0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;

     -- n8_MUX[uxn_opcodes_h_l2019_c7_3712] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2019_c7_3712_cond <= VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_cond;
     n8_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue;
     n8_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_return_output := n8_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2019_c7_3712] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2022_c7_0bd0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2019_c7_3712] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2022_c7_0bd0_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse := VAR_t8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2019_c7_3712] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2019_c7_3712] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2015_c7_e35b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2015_c7_e35b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;

     -- t8_MUX[uxn_opcodes_h_l2007_c2_cec3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond <= VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond;
     t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue;
     t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output := t8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2019_c7_3712] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_return_output := result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2019_c7_3712] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;

     -- n8_MUX[uxn_opcodes_h_l2015_c7_e35b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond <= VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_cond;
     n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue;
     n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output := n8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2019_c7_3712_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2012_c7_8196] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2015_c7_e35b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;

     -- n8_MUX[uxn_opcodes_h_l2012_c7_8196] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2012_c7_8196_cond <= VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_cond;
     n8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue;
     n8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output := n8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2012_c7_8196] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2015_c7_e35b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2015_c7_e35b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2015_c7_e35b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output := result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;

     -- Submodule level 5
     VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2015_c7_e35b_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l2007_c2_cec3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2012_c7_8196] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_return_output := result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2012_c7_8196] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2012_c7_8196] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l2007_c2_cec3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l2012_c7_8196] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;

     -- n8_MUX[uxn_opcodes_h_l2007_c2_cec3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond <= VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_cond;
     n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue;
     n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output := n8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;

     -- Submodule level 6
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l2012_c7_8196_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l2007_c2_cec3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l2007_c2_cec3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l2007_c2_cec3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output := result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l2007_c2_cec3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output;

     -- Submodule level 7
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2036_l2003_DUPLICATE_bab3 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2036_l2003_DUPLICATE_bab3_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_3345(
     result,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l2007_c2_cec3_return_output);

     -- Submodule level 8
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2036_l2003_DUPLICATE_bab3_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_3345_uxn_opcodes_h_l2036_l2003_DUPLICATE_bab3_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
