-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity lth_0CLK_226c8821 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end lth_0CLK_226c8821;
architecture arch of lth_0CLK_226c8821 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1906_c6_2f74]
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal n8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(7 downto 0);

-- result_is_ram_write_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
signal result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : signed(3 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(7 downto 0);

-- result_is_vram_write_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
signal result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1906_c2_55ea]
signal t8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1919_c11_fe8d]
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1919_c7_ec12]
signal n8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1919_c7_ec12]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1919_c7_ec12]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1919_c7_ec12]
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1919_c7_ec12]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1919_c7_ec12]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1919_c7_ec12]
signal t8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1922_c11_92ef]
signal BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1922_c7_aa15]
signal n8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1922_c7_aa15]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1922_c7_aa15]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1922_c7_aa15]
signal result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1922_c7_aa15]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1922_c7_aa15]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1922_c7_aa15]
signal t8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1925_c11_8f40]
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1925_c7_5c1c]
signal n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(7 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1925_c7_5c1c]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1925_c7_5c1c]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : signed(3 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1925_c7_5c1c]
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(7 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1925_c7_5c1c]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1925_c7_5c1c]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(0 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1927_c30_c08f]
signal sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_return_output : signed(3 downto 0);

-- BIN_OP_LT[uxn_opcodes_h_l1930_c21_b721]
signal BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_left : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_right : unsigned(7 downto 0);
signal BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1930_c21_0173]
signal MUX_uxn_opcodes_h_l1930_c21_0173_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1930_c21_0173_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1930_c21_0173_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1930_c21_0173_return_output : unsigned(7 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_a47b( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : signed;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.is_ram_write := ref_toks_1;
      base.is_opc_done := ref_toks_2;
      base.sp_relative_shift := ref_toks_3;
      base.is_stack_index_flipped := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.is_stack_write := ref_toks_6;
      base.is_pc_updated := ref_toks_7;
      base.u8_value := ref_toks_8;
      base.is_vram_write := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74
BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_left,
BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_right,
BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output);

-- n8_MUX_uxn_opcodes_h_l1906_c2_55ea
n8_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
n8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- t8_MUX_uxn_opcodes_h_l1906_c2_55ea
t8_MUX_uxn_opcodes_h_l1906_c2_55ea : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond,
t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue,
t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse,
t8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d
BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_left,
BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_right,
BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output);

-- n8_MUX_uxn_opcodes_h_l1919_c7_ec12
n8_MUX_uxn_opcodes_h_l1919_c7_ec12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond,
n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue,
n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse,
n8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_cond,
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output);

-- t8_MUX_uxn_opcodes_h_l1919_c7_ec12
t8_MUX_uxn_opcodes_h_l1919_c7_ec12 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond,
t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue,
t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse,
t8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef
BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_left,
BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_right,
BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output);

-- n8_MUX_uxn_opcodes_h_l1922_c7_aa15
n8_MUX_uxn_opcodes_h_l1922_c7_aa15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond,
n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue,
n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse,
n8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_cond,
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output);

-- t8_MUX_uxn_opcodes_h_l1922_c7_aa15
t8_MUX_uxn_opcodes_h_l1922_c7_aa15 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond,
t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue,
t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse,
t8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_left,
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_right,
BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output);

-- n8_MUX_uxn_opcodes_h_l1925_c7_5c1c
n8_MUX_uxn_opcodes_h_l1925_c7_5c1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond,
n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue,
n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse,
n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f
sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_ins,
sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_x,
sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_y,
sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_return_output);

-- BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721
BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721 : entity work.BIN_OP_LT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_left,
BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_right,
BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_return_output);

-- MUX_uxn_opcodes_h_l1930_c21_0173
MUX_uxn_opcodes_h_l1930_c21_0173 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1930_c21_0173_cond,
MUX_uxn_opcodes_h_l1930_c21_0173_iftrue,
MUX_uxn_opcodes_h_l1930_c21_0173_iffalse,
MUX_uxn_opcodes_h_l1930_c21_0173_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output,
 n8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 t8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output,
 n8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output,
 t8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output,
 n8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output,
 t8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output,
 n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output,
 sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_return_output,
 BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_return_output,
 MUX_uxn_opcodes_h_l1930_c21_0173_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1911_c3_b491 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1916_c3_5de0 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(0 downto 0);
 variable VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1920_c3_1152 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_4a87 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1930_c21_0173_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1930_c21_0173_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1930_c21_0173_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1930_c21_0173_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1925_l1919_l1922_DUPLICATE_bec0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_69db_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5d99_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5485_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_134b_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1934_l1902_DUPLICATE_3285_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_4a87 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1929_c3_4a87;
     VAR_MUX_uxn_opcodes_h_l1930_c21_0173_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_y := resize(to_signed(-1, 2), 4);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1911_c3_b491 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1911_c3_b491;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1916_c3_5de0 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1916_c3_5de0;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_right := to_unsigned(2, 2);
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_right := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1930_c21_0173_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_right := to_unsigned(3, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1920_c3_1152 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1920_c3_1152;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_left := VAR_phase;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1906_c6_2f74] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_left;
     BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output := BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5485 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5485_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1925_c11_8f40] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_left;
     BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output := BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_69db LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_69db_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1925_l1919_l1922_DUPLICATE_bec0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1925_l1919_l1922_DUPLICATE_bec0_return_output := result.u8_value;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_134b LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_134b_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1922_c11_92ef] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_left;
     BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output := BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output;

     -- result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output := result.is_pc_updated;

     -- result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output := result.is_stack_index_flipped;

     -- BIN_OP_LT[uxn_opcodes_h_l1930_c21_b721] LATENCY=0
     -- Inputs
     BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_left <= VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_left;
     BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_right <= VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_right;
     -- Outputs
     VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_return_output := BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_return_output;

     -- result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output := result.is_ram_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1919_c11_fe8d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_left;
     BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output := BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1927_c30_c08f] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_ins;
     sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_x;
     sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_return_output := sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5d99 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5d99_return_output := result.sp_relative_shift;

     -- result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output := result.is_vram_write;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1906_c6_2f74_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1919_c11_fe8d_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1922_c11_92ef_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1925_c11_8f40_return_output;
     VAR_MUX_uxn_opcodes_h_l1930_c21_0173_cond := VAR_BIN_OP_LT_uxn_opcodes_h_l1930_c21_b721_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5d99_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5d99_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5d99_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_69db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_69db_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_69db_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5485_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5485_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1925_l1919_l1922_DUPLICATE_5485_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_134b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1925_l1922_DUPLICATE_134b_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1925_l1919_l1922_DUPLICATE_bec0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1925_l1919_l1922_DUPLICATE_bec0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1925_l1919_l1922_DUPLICATE_bec0_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1906_l1925_l1919_l1922_DUPLICATE_bec0_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_is_pc_updated_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output;
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_is_ram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_ram_write_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_is_stack_index_flipped_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output;
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_is_vram_write_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_opcode_result_t_is_vram_write_d41d_uxn_opcodes_h_l1906_c2_55ea_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1927_c30_c08f_return_output;
     -- MUX[uxn_opcodes_h_l1930_c21_0173] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1930_c21_0173_cond <= VAR_MUX_uxn_opcodes_h_l1930_c21_0173_cond;
     MUX_uxn_opcodes_h_l1930_c21_0173_iftrue <= VAR_MUX_uxn_opcodes_h_l1930_c21_0173_iftrue;
     MUX_uxn_opcodes_h_l1930_c21_0173_iffalse <= VAR_MUX_uxn_opcodes_h_l1930_c21_0173_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1930_c21_0173_return_output := MUX_uxn_opcodes_h_l1930_c21_0173_return_output;

     -- t8_MUX[uxn_opcodes_h_l1922_c7_aa15] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond <= VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond;
     t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue;
     t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output := t8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;

     -- result_is_vram_write_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1925_c7_5c1c] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;

     -- result_is_ram_write_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- n8_MUX[uxn_opcodes_h_l1925_c7_5c1c] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond;
     n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue;
     n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output := n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1925_c7_5c1c] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1925_c7_5c1c] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1925_c7_5c1c] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue := VAR_MUX_uxn_opcodes_h_l1930_c21_0173_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1925_c7_5c1c] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output := result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1922_c7_aa15] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;

     -- t8_MUX[uxn_opcodes_h_l1919_c7_ec12] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond <= VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond;
     t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue;
     t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output := t8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1922_c7_aa15] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1922_c7_aa15] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1922_c7_aa15] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;

     -- n8_MUX[uxn_opcodes_h_l1922_c7_aa15] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond <= VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_cond;
     n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue;
     n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output := n8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1925_c7_5c1c_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1919_c7_ec12] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1922_c7_aa15] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output := result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1919_c7_ec12] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1919_c7_ec12] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;

     -- t8_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := t8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- n8_MUX[uxn_opcodes_h_l1919_c7_ec12] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond <= VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_cond;
     n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue;
     n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output := n8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1919_c7_ec12] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1922_c7_aa15_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;
     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- n8_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := n8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1919_c7_ec12] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output := result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1919_c7_ec12_return_output;
     -- result_u8_value_MUX[uxn_opcodes_h_l1906_c2_55ea] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output := result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1934_l1902_DUPLICATE_3285 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1934_l1902_DUPLICATE_3285_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_a47b(
     result,
     VAR_result_is_ram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output,
     VAR_result_is_vram_write_MUX_uxn_opcodes_h_l1906_c2_55ea_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1934_l1902_DUPLICATE_3285_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_a47b_uxn_opcodes_h_l1934_l1902_DUPLICATE_3285_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
