-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 39
entity gth_0CLK_7883ef49 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end gth_0CLK_7883ef49;
architecture arch of gth_0CLK_7883ef49 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1784_c6_9bcf]
signal BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1784_c2_123a]
signal n8_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1784_c2_123a]
signal result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1784_c2_123a]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1784_c2_123a]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1784_c2_123a]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1784_c2_123a]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1784_c2_123a]
signal t8_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1791_c11_9b84]
signal BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1791_c7_2a42]
signal n8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1791_c7_2a42]
signal result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1791_c7_2a42]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1791_c7_2a42]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1791_c7_2a42]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1791_c7_2a42]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1791_c7_2a42]
signal t8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1794_c11_eb96]
signal BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1794_c7_f9fa]
signal n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1794_c7_f9fa]
signal result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1794_c7_f9fa]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1794_c7_f9fa]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1794_c7_f9fa]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1794_c7_f9fa]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : signed(3 downto 0);

-- t8_MUX[uxn_opcodes_h_l1794_c7_f9fa]
signal t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1797_c11_e252]
signal BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1797_c7_c5ff]
signal n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1797_c7_c5ff]
signal result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(7 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1797_c7_c5ff]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1797_c7_c5ff]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1797_c7_c5ff]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1797_c7_c5ff]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1800_c30_7741]
signal sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_return_output : signed(3 downto 0);

-- BIN_OP_GT[uxn_opcodes_h_l1803_c21_19e9]
signal BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_left : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_right : unsigned(7 downto 0);
signal BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1803_c21_d75f]
signal MUX_uxn_opcodes_h_l1803_c21_d75f_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1803_c21_d75f_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1803_c21_d75f_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1803_c21_d75f_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1805_c11_34ee]
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1805_c7_3730]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1805_c7_3730]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1805_c7_3730]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_return_output : signed(3 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_eae7( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_stack_write := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.stack_address_sp_offset := ref_toks_4;
      base.sp_relative_shift := ref_toks_5;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf
BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_left,
BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_right,
BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output);

-- n8_MUX_uxn_opcodes_h_l1784_c2_123a
n8_MUX_uxn_opcodes_h_l1784_c2_123a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1784_c2_123a_cond,
n8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue,
n8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse,
n8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a
result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_cond,
result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a
result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a
result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a
result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_return_output);

-- t8_MUX_uxn_opcodes_h_l1784_c2_123a
t8_MUX_uxn_opcodes_h_l1784_c2_123a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1784_c2_123a_cond,
t8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue,
t8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse,
t8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84
BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84 : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_left,
BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_right,
BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output);

-- n8_MUX_uxn_opcodes_h_l1791_c7_2a42
n8_MUX_uxn_opcodes_h_l1791_c7_2a42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond,
n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue,
n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse,
n8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42
result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_cond,
result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42
result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42
result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42
result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output);

-- t8_MUX_uxn_opcodes_h_l1791_c7_2a42
t8_MUX_uxn_opcodes_h_l1791_c7_2a42 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond,
t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue,
t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse,
t8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96
BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_left,
BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_right,
BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output);

-- n8_MUX_uxn_opcodes_h_l1794_c7_f9fa
n8_MUX_uxn_opcodes_h_l1794_c7_f9fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond,
n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue,
n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse,
n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa
result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond,
result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa
result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa
result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa
result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output);

-- t8_MUX_uxn_opcodes_h_l1794_c7_f9fa
t8_MUX_uxn_opcodes_h_l1794_c7_f9fa : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond,
t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue,
t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse,
t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252
BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_left,
BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_right,
BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output);

-- n8_MUX_uxn_opcodes_h_l1797_c7_c5ff
n8_MUX_uxn_opcodes_h_l1797_c7_c5ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond,
n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue,
n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse,
n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff
result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond,
result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff
result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff
result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff
result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1800_c30_7741
sp_relative_shift_uxn_opcodes_h_l1800_c30_7741 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_ins,
sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_x,
sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_y,
sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_return_output);

-- BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9
BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9 : entity work.BIN_OP_GT_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_left,
BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_right,
BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_return_output);

-- MUX_uxn_opcodes_h_l1803_c21_d75f
MUX_uxn_opcodes_h_l1803_c21_d75f : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1803_c21_d75f_cond,
MUX_uxn_opcodes_h_l1803_c21_d75f_iftrue,
MUX_uxn_opcodes_h_l1803_c21_d75f_iffalse,
MUX_uxn_opcodes_h_l1803_c21_d75f_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_left,
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_right,
BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output,
 n8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
 t8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output,
 n8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output,
 t8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output,
 n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output,
 t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output,
 n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output,
 sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_return_output,
 BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_return_output,
 MUX_uxn_opcodes_h_l1803_c21_d75f_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1788_c3_cc25 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1792_c3_6fe4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_712e : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_iffalse : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l1806_c3_8229 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1784_l1797_l1791_l1794_DUPLICATE_225e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_a14b_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_b1ca_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1797_l1791_l1805_l1794_DUPLICATE_98f4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1797_l1794_DUPLICATE_8f0d_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1811_l1780_DUPLICATE_97b4_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_right := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1788_c3_cc25 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1788_c3_cc25;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1792_c3_6fe4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1792_c3_6fe4;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue := to_unsigned(1, 1);
     VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_iftrue := resize(to_unsigned(1, 1), 8);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l1806_c3_8229 := signed(std_logic_vector(resize(to_unsigned(0, 1), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l1806_c3_8229;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_right := to_unsigned(4, 3);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_right := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_712e := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1802_c3_712e;
     VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_iffalse := resize(to_unsigned(0, 1), 8);
     VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_y := resize(to_signed(-1, 2), 4);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_left := VAR_phase;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse := t8;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_a14b LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_a14b_return_output := result.is_stack_write;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1797_l1794_DUPLICATE_8f0d LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1797_l1794_DUPLICATE_8f0d_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1784_c6_9bcf] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_left;
     BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output := BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1784_l1797_l1791_l1794_DUPLICATE_225e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1784_l1797_l1791_l1794_DUPLICATE_225e_return_output := result.u8_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l1791_c11_9b84] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_left;
     BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output := BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_b1ca LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_b1ca_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1797_l1791_l1805_l1794_DUPLICATE_98f4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1797_l1791_l1805_l1794_DUPLICATE_98f4_return_output := result.is_opc_done;

     -- sp_relative_shift[uxn_opcodes_h_l1800_c30_7741] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_ins;
     sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_x;
     sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_return_output := sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1794_c11_eb96] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_left;
     BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output := BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output;

     -- BIN_OP_GT[uxn_opcodes_h_l1803_c21_19e9] LATENCY=0
     -- Inputs
     BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_left <= VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_left;
     BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_right <= VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_right;
     -- Outputs
     VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_return_output := BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1797_c11_e252] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_left;
     BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output := BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1805_c11_34ee] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_left;
     BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output := BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output;

     -- Submodule level 1
     VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1784_c6_9bcf_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1791_c11_9b84_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1794_c11_eb96_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1797_c11_e252_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1805_c11_34ee_return_output;
     VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_cond := VAR_BIN_OP_GT_uxn_opcodes_h_l1803_c21_19e9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_b1ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_b1ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_b1ca_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_b1ca_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1797_l1791_l1805_l1794_DUPLICATE_98f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1797_l1791_l1805_l1794_DUPLICATE_98f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1797_l1791_l1805_l1794_DUPLICATE_98f4_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1797_l1791_l1805_l1794_DUPLICATE_98f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_a14b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_a14b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_a14b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1784_l1791_l1805_l1794_DUPLICATE_a14b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1797_l1794_DUPLICATE_8f0d_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1797_l1794_DUPLICATE_8f0d_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1784_l1797_l1791_l1794_DUPLICATE_225e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1784_l1797_l1791_l1794_DUPLICATE_225e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1784_l1797_l1791_l1794_DUPLICATE_225e_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1784_l1797_l1791_l1794_DUPLICATE_225e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1800_c30_7741_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1805_c7_3730] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_return_output;

     -- t8_MUX[uxn_opcodes_h_l1794_c7_f9fa] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond <= VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond;
     t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue;
     t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output := t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;

     -- n8_MUX[uxn_opcodes_h_l1797_c7_c5ff] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond <= VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond;
     n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue;
     n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output := n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1805_c7_3730] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_return_output;

     -- MUX[uxn_opcodes_h_l1803_c21_d75f] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1803_c21_d75f_cond <= VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_cond;
     MUX_uxn_opcodes_h_l1803_c21_d75f_iftrue <= VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_iftrue;
     MUX_uxn_opcodes_h_l1803_c21_d75f_iffalse <= VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_return_output := MUX_uxn_opcodes_h_l1803_c21_d75f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1805_c7_3730] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1797_c7_c5ff] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue := VAR_MUX_uxn_opcodes_h_l1803_c21_d75f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1805_c7_3730_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1805_c7_3730_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1805_c7_3730_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1797_c7_c5ff] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1797_c7_c5ff] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1797_c7_c5ff] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output := result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;

     -- t8_MUX[uxn_opcodes_h_l1791_c7_2a42] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond <= VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond;
     t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue;
     t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output := t8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1797_c7_c5ff] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1794_c7_f9fa] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;

     -- n8_MUX[uxn_opcodes_h_l1794_c7_f9fa] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond <= VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond;
     n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue;
     n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output := n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1797_c7_c5ff_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1794_c7_f9fa] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1794_c7_f9fa] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output := result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;

     -- t8_MUX[uxn_opcodes_h_l1784_c2_123a] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1784_c2_123a_cond <= VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_cond;
     t8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue;
     t8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output := t8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;

     -- n8_MUX[uxn_opcodes_h_l1791_c7_2a42] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond <= VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_cond;
     n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue;
     n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output := n8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1791_c7_2a42] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1794_c7_f9fa] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1794_c7_f9fa] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1794_c7_f9fa_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;
     -- result_is_opc_done_MUX[uxn_opcodes_h_l1791_c7_2a42] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1791_c7_2a42] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1791_c7_2a42] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;

     -- n8_MUX[uxn_opcodes_h_l1784_c2_123a] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1784_c2_123a_cond <= VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_cond;
     n8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue;
     n8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output := n8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1791_c7_2a42] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output := result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1784_c2_123a] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1791_c7_2a42_return_output;
     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1784_c2_123a] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1784_c2_123a] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_return_output := result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1784_c2_123a] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1784_c2_123a] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1811_l1780_DUPLICATE_97b4 LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1811_l1780_DUPLICATE_97b4_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_eae7(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1784_c2_123a_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1784_c2_123a_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1811_l1780_DUPLICATE_97b4_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_eae7_uxn_opcodes_h_l1811_l1780_DUPLICATE_97b4_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
