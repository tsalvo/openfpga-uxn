-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 47
entity jsr2_0CLK_fedec265 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 pc : in unsigned(15 downto 0);
 previous_stack_read : in unsigned(15 downto 0);
 return_output : out opcode_result_t);
end jsr2_0CLK_fedec265;
architecture arch of jsr2_0CLK_fedec265 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t16 : unsigned(15 downto 0) := to_unsigned(0, 16);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t16 : unsigned(15 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l741_c6_86cd]
signal BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l741_c2_e584]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l741_c2_e584]
signal t16_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l749_c11_1d8e]
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l749_c7_434f]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l749_c7_434f]
signal t16_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(15 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l751_c30_edf5]
signal sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l753_c11_4de3]
signal BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(15 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : signed(3 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(3 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l753_c7_32d3]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);

-- t16_MUX[uxn_opcodes_h_l753_c7_32d3]
signal t16_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
signal t16_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(15 downto 0);
signal t16_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(15 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l761_c11_d4ae]
signal BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l761_c7_36c9]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);

-- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l761_c7_36c9]
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);

-- result_u16_value_MUX[uxn_opcodes_h_l761_c7_36c9]
signal result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(15 downto 0);
signal result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(15 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l761_c7_36c9]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l761_c7_36c9]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l761_c7_36c9]
signal result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l761_c7_36c9]
signal result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l768_c11_2b57]
signal BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output : unsigned(0 downto 0);

-- result_is_pc_updated_MUX[uxn_opcodes_h_l768_c7_de83]
signal result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_cond : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iftrue : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iffalse : unsigned(0 downto 0);
signal result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l768_c7_de83]
signal result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_return_output : unsigned(0 downto 0);

-- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l768_c7_de83]
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_cond : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iftrue : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iffalse : unsigned(0 downto 0);
signal result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_4b08( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : signed;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u16_value := ref_toks_1;
      base.is_pc_updated := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.sp_relative_shift := ref_toks_4;
      base.is_stack_write := ref_toks_5;
      base.stack_address_sp_offset := ref_toks_6;
      base.is_sp_shift := ref_toks_7;
      base.is_stack_index_flipped := ref_toks_8;
      base.is_stack_operation_16bit := ref_toks_9;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd
BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_left,
BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_right,
BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584
result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584
result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584
result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584
result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584
result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584
result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- t16_MUX_uxn_opcodes_h_l741_c2_e584
t16_MUX_uxn_opcodes_h_l741_c2_e584 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l741_c2_e584_cond,
t16_MUX_uxn_opcodes_h_l741_c2_e584_iftrue,
t16_MUX_uxn_opcodes_h_l741_c2_e584_iffalse,
t16_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e
BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_left,
BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_right,
BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f
result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f
result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- t16_MUX_uxn_opcodes_h_l749_c7_434f
t16_MUX_uxn_opcodes_h_l749_c7_434f : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l749_c7_434f_cond,
t16_MUX_uxn_opcodes_h_l749_c7_434f_iftrue,
t16_MUX_uxn_opcodes_h_l749_c7_434f_iffalse,
t16_MUX_uxn_opcodes_h_l749_c7_434f_return_output);

-- sp_relative_shift_uxn_opcodes_h_l751_c30_edf5
sp_relative_shift_uxn_opcodes_h_l751_c30_edf5 : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_ins,
sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_x,
sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_y,
sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3
BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_left,
BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_right,
BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3
result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3
result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3
result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3
result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3
result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3
result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- t16_MUX_uxn_opcodes_h_l753_c7_32d3
t16_MUX_uxn_opcodes_h_l753_c7_32d3 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
t16_MUX_uxn_opcodes_h_l753_c7_32d3_cond,
t16_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue,
t16_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse,
t16_MUX_uxn_opcodes_h_l753_c7_32d3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae
BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_left,
BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_right,
BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9
result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_return_output);

-- result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_cond,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse,
result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_return_output);

-- result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9
result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9 : entity work.MUX_uint1_t_uint16_t_uint16_t_0CLK_de264c78 port map (
result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_cond,
result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue,
result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse,
result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9
result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9
result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9
result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57
BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_left,
BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_right,
BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output);

-- result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83
result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_cond,
result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iftrue,
result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iffalse,
result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83
result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_return_output);

-- result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_cond,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iftrue,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iffalse,
result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 pc,
 previous_stack_read,
 -- Registers
 t16,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 t16_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 t16_MUX_uxn_opcodes_h_l749_c7_434f_return_output,
 sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 t16_MUX_uxn_opcodes_h_l753_c7_32d3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_return_output,
 result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_return_output,
 result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output,
 result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_return_output,
 result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_pc : unsigned(15 downto 0);
 variable VAR_previous_stack_read : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l746_c3_4dd5 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_return_output : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_return_output : signed(3 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_uxn_opcodes_h_l756_c3_1a93 : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l758_c3_d163 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse : unsigned(15 downto 0);
 variable VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(15 downto 0);
 variable VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_edce_return_output : unsigned(15 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l749_l768_l753_l741_DUPLICATE_4c56_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l753_l741_DUPLICATE_ea47_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_9a88_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l761_l753_l741_DUPLICATE_66cb_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l761_l749_l768_l741_DUPLICATE_3e17_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l761_l749_l768_l753_DUPLICATE_62ef_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l749_l753_DUPLICATE_444a_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l761_l749_l753_DUPLICATE_18c2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l737_l774_DUPLICATE_c29c_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t16 : unsigned(15 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t16 := t16;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_right := to_unsigned(1, 1);
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_right := to_unsigned(3, 2);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := to_unsigned(1, 1);
     VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_y := resize(to_signed(-2, 3), 4);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iftrue := to_unsigned(0, 1);
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := to_unsigned(1, 1);
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue := to_unsigned(0, 1);
     VAR_result_sp_relative_shift_uxn_opcodes_h_l756_c3_1a93 := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := VAR_result_sp_relative_shift_uxn_opcodes_h_l756_c3_1a93;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l758_c3_d163 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l758_c3_d163;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue := to_unsigned(0, 1);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_right := to_unsigned(2, 2);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l746_c3_4dd5 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l746_c3_4dd5;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_right := to_unsigned(4, 3);
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_right := to_unsigned(0, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue := to_unsigned(0, 1);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_pc := pc;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_ins := VAR_ins;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := VAR_pc;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_left := VAR_phase;
     VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := VAR_previous_stack_read;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := t16;
     VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := t16;
     -- CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l749_l768_l753_l741_DUPLICATE_4c56 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l749_l768_l753_l741_DUPLICATE_4c56_return_output := result.is_pc_updated;

     -- sp_relative_shift[uxn_opcodes_h_l751_c30_edf5] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_ins;
     sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_x <= VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_x;
     sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_y <= VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_return_output := sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l761_c11_d4ae] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_left;
     BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output := BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l768_c11_2b57] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_left;
     BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output := BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l761_l753_l741_DUPLICATE_66cb LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l761_l753_l741_DUPLICATE_66cb_return_output := result.is_sp_shift;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l761_l749_l753_DUPLICATE_18c2 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l761_l749_l753_DUPLICATE_18c2_return_output := result.is_stack_operation_16bit;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_9a88 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_9a88_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l749_c11_1d8e] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_left;
     BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output := BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l761_l749_l768_l753_DUPLICATE_62ef LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l761_l749_l768_l753_DUPLICATE_62ef_return_output := result.is_opc_done;

     -- BIN_OP_EQ[uxn_opcodes_h_l753_c11_4de3] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_left;
     BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output := BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l749_l753_DUPLICATE_444a LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l749_l753_DUPLICATE_444a_return_output := result.stack_address_sp_offset;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l761_l749_l768_l741_DUPLICATE_3e17 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l761_l749_l768_l741_DUPLICATE_3e17_return_output := result.is_stack_index_flipped;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l753_l741_DUPLICATE_ea47 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l753_l741_DUPLICATE_ea47_return_output := result.sp_relative_shift;

     -- CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_edce LATENCY=0
     VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_edce_return_output := result.u16_value;

     -- BIN_OP_EQ[uxn_opcodes_h_l741_c6_86cd] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_left;
     BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output := BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;

     -- Submodule level 1
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l741_c6_86cd_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l749_c11_1d8e_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l753_c11_4de3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l761_c11_d4ae_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l768_c11_2b57_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l753_l741_DUPLICATE_ea47_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l753_l741_DUPLICATE_ea47_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_edce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_edce_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse := VAR_CONST_REF_RD_uint16_t_opcode_result_t_u16_value_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_edce_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l761_l749_l768_l753_DUPLICATE_62ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l761_l749_l768_l753_DUPLICATE_62ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l761_l749_l768_l753_DUPLICATE_62ef_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l761_l749_l768_l753_DUPLICATE_62ef_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l749_l768_l753_l741_DUPLICATE_4c56_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l749_l768_l753_l741_DUPLICATE_4c56_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l749_l768_l753_l741_DUPLICATE_4c56_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_pc_updated_d41d_uxn_opcodes_h_l749_l768_l753_l741_DUPLICATE_4c56_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l761_l753_l741_DUPLICATE_66cb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l761_l753_l741_DUPLICATE_66cb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l761_l753_l741_DUPLICATE_66cb_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l761_l749_l768_l741_DUPLICATE_3e17_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l761_l749_l768_l741_DUPLICATE_3e17_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l761_l749_l768_l741_DUPLICATE_3e17_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_index_flipped_d41d_uxn_opcodes_h_l761_l749_l768_l741_DUPLICATE_3e17_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l761_l749_l753_DUPLICATE_18c2_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l761_l749_l753_DUPLICATE_18c2_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_operation_16bit_d41d_uxn_opcodes_h_l761_l749_l753_DUPLICATE_18c2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_9a88_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_9a88_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l761_l749_l741_DUPLICATE_9a88_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l749_l753_DUPLICATE_444a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l749_l753_DUPLICATE_444a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l751_c30_edf5_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l761_c7_36c9] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l761_c7_36c9] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l768_c7_de83] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l761_c7_36c9] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l761_c7_36c9] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_cond;
     result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_return_output := result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l768_c7_de83] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l768_c7_de83] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_return_output;

     -- t16_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     t16_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     t16_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := t16_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- Submodule level 2
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l768_c7_de83_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l768_c7_de83_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l768_c7_de83_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_t16_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l761_c7_36c9] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l761_c7_36c9] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l761_c7_36c9] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- t16_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     t16_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     t16_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_return_output := t16_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- Submodule level 3
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l761_c7_36c9_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_t16_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     -- result_u16_value_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- t16_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     t16_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     t16_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     t16_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_return_output := t16_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l753_c7_32d3] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- Submodule level 4
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l753_c7_32d3_return_output;
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_u16_value_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     REG_VAR_t16 := VAR_t16_MUX_uxn_opcodes_h_l741_c2_e584_return_output;
     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- result_is_pc_updated_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l749_c7_434f] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_return_output;

     -- result_is_stack_operation_16bit_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- result_u16_value_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- Submodule level 5
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iffalse := VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l749_c7_434f_return_output;
     -- result_is_pc_updated_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- result_is_stack_index_flipped_MUX[uxn_opcodes_h_l741_c2_e584] LATENCY=0
     -- Inputs
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_cond <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_cond;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iftrue <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iftrue;
     result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iffalse <= VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_iffalse;
     -- Outputs
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_return_output := result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l737_l774_DUPLICATE_c29c LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l737_l774_DUPLICATE_c29c_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_4b08(
     result,
     VAR_result_u16_value_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
     VAR_result_is_pc_updated_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
     VAR_result_is_stack_index_flipped_MUX_uxn_opcodes_h_l741_c2_e584_return_output,
     VAR_result_is_stack_operation_16bit_MUX_uxn_opcodes_h_l741_c2_e584_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l737_l774_DUPLICATE_c29c_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_4b08_uxn_opcodes_h_l737_l774_DUPLICATE_c29c_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t16 <= REG_VAR_t16;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t16 <= REG_COMB_t16;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
