-- Timing params:
--   Fixed?: True
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 45
entity neq_0CLK_85d5529e is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 phase : in unsigned(7 downto 0);
 ins : in unsigned(7 downto 0);
 previous_stack_read : in unsigned(7 downto 0);
 return_output : out opcode_result_t);
end neq_0CLK_85d5529e;
architecture arch of neq_0CLK_85d5529e is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal t8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal n8 : unsigned(7 downto 0) := to_unsigned(0, 8);
signal result : opcode_result_t := opcode_result_t_NULL;
signal REG_COMB_t8 : unsigned(7 downto 0);
signal REG_COMB_n8 : unsigned(7 downto 0);
signal REG_COMB_result : opcode_result_t;

-- Each function instance gets signals
-- BIN_OP_EQ[uxn_opcodes_h_l1188_c6_088f]
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1188_c1_d3da]
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1188_c2_1fd0]
signal t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1188_c2_1fd0]
signal n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1188_c2_1fd0]
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1188_c2_1fd0]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1188_c2_1fd0]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1188_c2_1fd0]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1188_c2_1fd0]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1188_c2_1fd0]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : signed(3 downto 0);

-- printf_uxn_opcodes_h_l1189_c3_cace[uxn_opcodes_h_l1189_c3_cace]
signal printf_uxn_opcodes_h_l1189_c3_cace_uxn_opcodes_h_l1189_c3_cace_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1193_c11_300a]
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_right : unsigned(0 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1193_c7_b9eb]
signal t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1193_c7_b9eb]
signal n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1193_c7_b9eb]
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1193_c7_b9eb]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1193_c7_b9eb]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1193_c7_b9eb]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1193_c7_b9eb]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1193_c7_b9eb]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1196_c11_7639]
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output : unsigned(0 downto 0);

-- t8_MUX[uxn_opcodes_h_l1196_c7_17d3]
signal t8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(7 downto 0);
signal t8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(7 downto 0);

-- n8_MUX[uxn_opcodes_h_l1196_c7_17d3]
signal n8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1196_c7_17d3]
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1196_c7_17d3]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1196_c7_17d3]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1196_c7_17d3]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1196_c7_17d3]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1196_c7_17d3]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_e9e2]
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_right : unsigned(1 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output : unsigned(0 downto 0);

-- n8_MUX[uxn_opcodes_h_l1199_c7_147b]
signal n8_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(7 downto 0);
signal n8_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(7 downto 0);

-- result_u8_value_MUX[uxn_opcodes_h_l1199_c7_147b]
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(7 downto 0);
signal result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(7 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1199_c7_147b]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_147b]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_147b]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(0 downto 0);

-- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1199_c7_147b]
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(3 downto 0);
signal result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(3 downto 0);

-- result_sp_relative_shift_MUX[uxn_opcodes_h_l1199_c7_147b]
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : signed(3 downto 0);
signal result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : signed(3 downto 0);

-- sp_relative_shift[uxn_opcodes_h_l1202_c30_cd7c]
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_ins : unsigned(7 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_x : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_y : signed(3 downto 0);
signal sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_return_output : signed(3 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1205_c21_6d46]
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_right : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_return_output : unsigned(0 downto 0);

-- MUX[uxn_opcodes_h_l1205_c21_cd39]
signal MUX_uxn_opcodes_h_l1205_c21_cd39_cond : unsigned(0 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_cd39_iftrue : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_cd39_iffalse : unsigned(7 downto 0);
signal MUX_uxn_opcodes_h_l1205_c21_cd39_return_output : unsigned(7 downto 0);

-- BIN_OP_EQ[uxn_opcodes_h_l1207_c11_17d6]
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_left : unsigned(7 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_right : unsigned(2 downto 0);
signal BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output : unsigned(0 downto 0);

-- result_is_sp_shift_MUX[uxn_opcodes_h_l1207_c7_b9d2]
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse : unsigned(0 downto 0);
signal result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output : unsigned(0 downto 0);

-- result_is_opc_done_MUX[uxn_opcodes_h_l1207_c7_b9d2]
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse : unsigned(0 downto 0);
signal result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output : unsigned(0 downto 0);

-- result_is_stack_write_MUX[uxn_opcodes_h_l1207_c7_b9d2]
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse : unsigned(0 downto 0);
signal result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output : unsigned(0 downto 0);

function CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2( ref_toks_0 : opcode_result_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : signed) return opcode_result_t is
 
  variable base : opcode_result_t; 
  variable return_output : opcode_result_t;
begin
      base := ref_toks_0;
      base.u8_value := ref_toks_1;
      base.is_sp_shift := ref_toks_2;
      base.is_opc_done := ref_toks_3;
      base.is_stack_write := ref_toks_4;
      base.stack_address_sp_offset := ref_toks_5;
      base.sp_relative_shift := ref_toks_6;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_left,
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_right,
BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output);

-- TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_cond,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iftrue,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iffalse,
TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_return_output);

-- t8_MUX_uxn_opcodes_h_l1188_c2_1fd0
t8_MUX_uxn_opcodes_h_l1188_c2_1fd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond,
t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue,
t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse,
t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

-- n8_MUX_uxn_opcodes_h_l1188_c2_1fd0
n8_MUX_uxn_opcodes_h_l1188_c2_1fd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond,
n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue,
n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse,
n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

-- printf_uxn_opcodes_h_l1189_c3_cace_uxn_opcodes_h_l1189_c3_cace
printf_uxn_opcodes_h_l1189_c3_cace_uxn_opcodes_h_l1189_c3_cace : entity work.printf_uxn_opcodes_h_l1189_c3_cace_0CLK_de264c78 port map (
printf_uxn_opcodes_h_l1189_c3_cace_uxn_opcodes_h_l1189_c3_cace_CLOCK_ENABLE);

-- BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a : entity work.BIN_OP_EQ_uint8_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_left,
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_right,
BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output);

-- t8_MUX_uxn_opcodes_h_l1193_c7_b9eb
t8_MUX_uxn_opcodes_h_l1193_c7_b9eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond,
t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue,
t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse,
t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output);

-- n8_MUX_uxn_opcodes_h_l1193_c7_b9eb
n8_MUX_uxn_opcodes_h_l1193_c7_b9eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond,
n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue,
n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse,
n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_left,
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_right,
BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output);

-- t8_MUX_uxn_opcodes_h_l1196_c7_17d3
t8_MUX_uxn_opcodes_h_l1196_c7_17d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
t8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond,
t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue,
t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse,
t8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output);

-- n8_MUX_uxn_opcodes_h_l1196_c7_17d3
n8_MUX_uxn_opcodes_h_l1196_c7_17d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond,
n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue,
n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse,
n8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_cond,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3 : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3 : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2 : entity work.BIN_OP_EQ_uint8_t_uint2_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_left,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_right,
BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output);

-- n8_MUX_uxn_opcodes_h_l1199_c7_147b
n8_MUX_uxn_opcodes_h_l1199_c7_147b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
n8_MUX_uxn_opcodes_h_l1199_c7_147b_cond,
n8_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue,
n8_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse,
n8_MUX_uxn_opcodes_h_l1199_c7_147b_return_output);

-- result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_cond,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse,
result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_return_output);

-- result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b : entity work.MUX_uint1_t_uint4_t_uint4_t_0CLK_de264c78 port map (
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_cond,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse,
result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_return_output);

-- result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b : entity work.MUX_uint1_t_int4_t_int4_t_0CLK_de264c78 port map (
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse,
result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output);

-- sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c
sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c : entity work.sp_relative_shift_0CLK_6f2c5aad port map (
sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_ins,
sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_x,
sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_y,
sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46 : entity work.BIN_OP_EQ_uint8_t_uint8_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_left,
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_right,
BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_return_output);

-- MUX_uxn_opcodes_h_l1205_c21_cd39
MUX_uxn_opcodes_h_l1205_c21_cd39 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
MUX_uxn_opcodes_h_l1205_c21_cd39_cond,
MUX_uxn_opcodes_h_l1205_c21_cd39_iftrue,
MUX_uxn_opcodes_h_l1205_c21_cd39_iffalse,
MUX_uxn_opcodes_h_l1205_c21_cd39_return_output);

-- BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6 : entity work.BIN_OP_EQ_uint8_t_uint3_t_0CLK_de264c78 port map (
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_left,
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_right,
BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output);

-- result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse,
result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output);

-- result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse,
result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output);

-- result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse,
result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output);



-- Combinatorial process for pipeline stages
process (
 CLOCK_ENABLE,
 -- Inputs
 phase,
 ins,
 previous_stack_read,
 -- Registers
 t8,
 n8,
 result,
 -- All submodule outputs
 BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output,
 TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_return_output,
 t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
 n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output,
 t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output,
 n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output,
 t8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output,
 n8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output,
 n8_MUX_uxn_opcodes_h_l1199_c7_147b_return_output,
 result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_return_output,
 result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_return_output,
 result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output,
 sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_return_output,
 MUX_uxn_opcodes_h_l1205_c21_cd39_return_output,
 BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output,
 result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output,
 result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output,
 result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : opcode_result_t;
 variable VAR_phase : unsigned(7 downto 0);
 variable VAR_ins : unsigned(7 downto 0);
 variable VAR_previous_stack_read : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iffalse : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_89f8 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond : unsigned(0 downto 0);
 variable VAR_printf_uxn_opcodes_h_l1189_c3_cace_uxn_opcodes_h_l1189_c3_cace_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_8de4 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output : unsigned(0 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(7 downto 0);
 variable VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output : unsigned(0 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(7 downto 0);
 variable VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(7 downto 0);
 variable VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_8d05 : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : unsigned(3 downto 0);
 variable VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse : signed(3 downto 0);
 variable VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond : unsigned(0 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_ins : unsigned(7 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_x : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_y : signed(3 downto 0);
 variable VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_return_output : signed(3 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_cond : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_iftrue : unsigned(7 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_iffalse : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_right : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_return_output : unsigned(0 downto 0);
 variable VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_left : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_right : unsigned(2 downto 0);
 variable VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse : unsigned(0 downto 0);
 variable VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_5112_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_11f4_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_b448_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_e580_return_output : signed(3 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_9ad9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_6790_return_output : unsigned(3 downto 0);
 variable VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1213_l1184_DUPLICATE_f02f_return_output : opcode_result_t;
 -- State registers comb logic variables
variable REG_VAR_t8 : unsigned(7 downto 0);
variable REG_VAR_n8 : unsigned(7 downto 0);
variable REG_VAR_result : opcode_result_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_t8 := t8;
  REG_VAR_n8 := n8;
  REG_VAR_result := result;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_right := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_8de4 := resize(to_unsigned(2, 2), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1194_c3_8de4;
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_8d05 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1204_c3_8d05;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue := to_unsigned(0, 1);
     VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_iffalse := resize(to_unsigned(1, 1), 8);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_right := to_unsigned(3, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_y := resize(to_signed(-1, 2), 4);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_right := to_unsigned(2, 2);
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_x := signed(std_logic_vector(resize(to_unsigned(2, 2), 4)));
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iffalse := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue := to_unsigned(0, 1);
     VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_89f8 := resize(to_unsigned(1, 1), 4);
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue := VAR_result_stack_address_sp_offset_uxn_opcodes_h_l1190_c3_89f8;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue := to_unsigned(1, 1);
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue := to_unsigned(0, 1);
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_right := to_unsigned(4, 3);
     VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_iftrue := resize(to_unsigned(0, 1), 8);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE := CLOCK_ENABLE;
     -- Mux in inputs
     VAR_phase := phase;
     VAR_ins := ins;
     VAR_previous_stack_read := previous_stack_read;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iftrue := VAR_CLOCK_ENABLE;
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_ins := VAR_ins;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue := n8;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse := n8;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_left := VAR_phase;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_left := VAR_previous_stack_read;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue := VAR_previous_stack_read;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue := VAR_previous_stack_read;
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_right := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue := t8;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse := t8;
     -- BIN_OP_EQ[uxn_opcodes_h_l1207_c11_17d6] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_left;
     BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output := BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1199_c11_e9e2] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_left;
     BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output := BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output;

     -- sp_relative_shift[uxn_opcodes_h_l1202_c30_cd7c] LATENCY=0
     -- Inputs
     sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_ins <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_ins;
     sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_x <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_x;
     sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_y <= VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_y;
     -- Outputs
     VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_return_output := sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_return_output;

     -- CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_6790 LATENCY=0
     VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_6790_return_output := result.stack_address_sp_offset;

     -- BIN_OP_EQ[uxn_opcodes_h_l1193_c11_300a] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_left;
     BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output := BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_11f4 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_11f4_return_output := result.is_sp_shift;

     -- CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_e580 LATENCY=0
     VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_e580_return_output := result.sp_relative_shift;

     -- BIN_OP_EQ[uxn_opcodes_h_l1188_c6_088f] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_left;
     BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output := BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;

     -- BIN_OP_EQ[uxn_opcodes_h_l1196_c11_7639] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_left;
     BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output := BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_b448 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_b448_return_output := result.is_stack_write;

     -- BIN_OP_EQ[uxn_opcodes_h_l1205_c21_6d46] LATENCY=0
     -- Inputs
     BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_left <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_left;
     BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_right <= VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_right;
     -- Outputs
     VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_return_output := BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_return_output;

     -- CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_9ad9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_9ad9_return_output := result.is_opc_done;

     -- CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_5112 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_5112_return_output := result.u8_value;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1188_c6_088f_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1193_c11_300a_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1196_c11_7639_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1199_c11_e9e2_return_output;
     VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1205_c21_6d46_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond := VAR_BIN_OP_EQ_uxn_opcodes_h_l1207_c11_17d6_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_e580_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_e580_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_e580_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse := VAR_CONST_REF_RD_int4_t_opcode_result_t_sp_relative_shift_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_e580_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_9ad9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_9ad9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_9ad9_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_opc_done_d41d_uxn_opcodes_h_l1199_l1193_l1207_l1196_DUPLICATE_9ad9_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_11f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_11f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_11f4_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_sp_shift_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_11f4_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_b448_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_b448_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_b448_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse := VAR_CONST_REF_RD_uint1_t_opcode_result_t_is_stack_write_d41d_uxn_opcodes_h_l1193_l1207_l1196_l1188_DUPLICATE_b448_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_6790_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse := VAR_CONST_REF_RD_uint4_t_opcode_result_t_stack_address_sp_offset_d41d_uxn_opcodes_h_l1199_l1196_DUPLICATE_6790_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_5112_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_5112_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_5112_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse := VAR_CONST_REF_RD_uint8_t_opcode_result_t_u8_value_d41d_uxn_opcodes_h_l1199_l1193_l1196_l1188_DUPLICATE_5112_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue := VAR_sp_relative_shift_uxn_opcodes_h_l1202_c30_cd7c_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1207_c7_b9d2] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1199_c7_147b] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1207_c7_b9d2] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1207_c7_b9d2] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output;

     -- MUX[uxn_opcodes_h_l1205_c21_cd39] LATENCY=0
     -- Inputs
     MUX_uxn_opcodes_h_l1205_c21_cd39_cond <= VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_cond;
     MUX_uxn_opcodes_h_l1205_c21_cd39_iftrue <= VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_iftrue;
     MUX_uxn_opcodes_h_l1205_c21_cd39_iffalse <= VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_iffalse;
     -- Outputs
     VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_return_output := MUX_uxn_opcodes_h_l1205_c21_cd39_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1199_c7_147b] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;

     -- t8_MUX[uxn_opcodes_h_l1196_c7_17d3] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond;
     t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue;
     t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output := t8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;

     -- n8_MUX[uxn_opcodes_h_l1199_c7_147b] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1199_c7_147b_cond <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_cond;
     n8_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue;
     n8_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_return_output := n8_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[uxn_opcodes_h_l1188_c1_d3da] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_cond;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iftrue;
     TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_return_output := TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_return_output;

     -- Submodule level 2
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue := VAR_MUX_uxn_opcodes_h_l1205_c21_cd39_return_output;
     VAR_printf_uxn_opcodes_h_l1189_c3_cace_uxn_opcodes_h_l1189_c3_cace_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_uxn_opcodes_h_l1188_c1_d3da_return_output;
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1207_c7_b9d2_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;
     -- n8_MUX[uxn_opcodes_h_l1196_c7_17d3] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_cond;
     n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue;
     n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output := n8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1199_c7_147b] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1199_c7_147b] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1199_c7_147b] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1199_c7_147b] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_return_output := result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1196_c7_17d3] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;

     -- t8_MUX[uxn_opcodes_h_l1193_c7_b9eb] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond;
     t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue;
     t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output := t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1196_c7_17d3] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;

     -- printf_uxn_opcodes_h_l1189_c3_cace[uxn_opcodes_h_l1189_c3_cace] LATENCY=0
     -- Clock enable
     printf_uxn_opcodes_h_l1189_c3_cace_uxn_opcodes_h_l1189_c3_cace_CLOCK_ENABLE <= VAR_printf_uxn_opcodes_h_l1189_c3_cace_uxn_opcodes_h_l1189_c3_cace_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- Submodule level 3
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1199_c7_147b_return_output;
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse := VAR_t8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1196_c7_17d3] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1196_c7_17d3] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1196_c7_17d3] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1196_c7_17d3] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output := result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1193_c7_b9eb] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;

     -- n8_MUX[uxn_opcodes_h_l1193_c7_b9eb] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond;
     n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue;
     n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output := n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;

     -- t8_MUX[uxn_opcodes_h_l1188_c2_1fd0] LATENCY=0
     -- Inputs
     t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond;
     t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue;
     t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse <= VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse;
     -- Outputs
     VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output := t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1193_c7_b9eb] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;

     -- Submodule level 4
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse := VAR_n8_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse := VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse := VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1196_c7_17d3_return_output;
     REG_VAR_t8 := VAR_t8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;
     -- result_is_stack_write_MUX[uxn_opcodes_h_l1193_c7_b9eb] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;

     -- result_stack_address_sp_offset_MUX[uxn_opcodes_h_l1188_c2_1fd0] LATENCY=0
     -- Inputs
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue;
     result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse <= VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse;
     -- Outputs
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output := result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;

     -- n8_MUX[uxn_opcodes_h_l1188_c2_1fd0] LATENCY=0
     -- Inputs
     n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond;
     n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue;
     n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse <= VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse;
     -- Outputs
     VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output := n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;

     -- result_sp_relative_shift_MUX[uxn_opcodes_h_l1188_c2_1fd0] LATENCY=0
     -- Inputs
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue;
     result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse <= VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse;
     -- Outputs
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output := result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1193_c7_b9eb] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output := result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1193_c7_b9eb] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;

     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1193_c7_b9eb] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;

     -- Submodule level 5
     REG_VAR_n8 := VAR_n8_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse := VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse := VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse := VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse := VAR_result_u8_value_MUX_uxn_opcodes_h_l1193_c7_b9eb_return_output;
     -- result_is_sp_shift_MUX[uxn_opcodes_h_l1188_c2_1fd0] LATENCY=0
     -- Inputs
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue;
     result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse <= VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse;
     -- Outputs
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output := result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;

     -- result_u8_value_MUX[uxn_opcodes_h_l1188_c2_1fd0] LATENCY=0
     -- Inputs
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond;
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue;
     result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse <= VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse;
     -- Outputs
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output := result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;

     -- result_is_stack_write_MUX[uxn_opcodes_h_l1188_c2_1fd0] LATENCY=0
     -- Inputs
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond;
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue;
     result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse <= VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse;
     -- Outputs
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output := result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;

     -- result_is_opc_done_MUX[uxn_opcodes_h_l1188_c2_1fd0] LATENCY=0
     -- Inputs
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_cond;
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iftrue;
     result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse <= VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_iffalse;
     -- Outputs
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output := result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output;

     -- Submodule level 6
     -- CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1213_l1184_DUPLICATE_f02f LATENCY=0
     VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1213_l1184_DUPLICATE_f02f_return_output := CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2(
     result,
     VAR_result_u8_value_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
     VAR_result_is_sp_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
     VAR_result_is_opc_done_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
     VAR_result_is_stack_write_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
     VAR_result_stack_address_sp_offset_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output,
     VAR_result_sp_relative_shift_MUX_uxn_opcodes_h_l1188_c2_1fd0_return_output);

     -- Submodule level 7
     REG_VAR_result := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1213_l1184_DUPLICATE_f02f_return_output;
     VAR_return_output := VAR_CONST_REF_RD_opcode_result_t_opcode_result_t_5cd2_uxn_opcodes_h_l1213_l1184_DUPLICATE_f02f_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_t8 <= REG_VAR_t8;
REG_COMB_n8 <= REG_VAR_n8;
REG_COMB_result <= REG_VAR_result;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if CLOCK_ENABLE(0)='1' then
     t8 <= REG_COMB_t8;
     n8 <= REG_COMB_n8;
     result <= REG_COMB_result;
 end if;
 end if;
end process;

end arch;
